module level_1(x, y, value);
    input [5:0] x;
    input [4:0] y;
    output [2:0] value;

    reg [2:0] value;
    always @(*)
    case (x)
        6'd0: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd7;
                5'd2: value = 3'd7;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd1: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd4;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd2: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd4;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd4;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd3: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd7;
                5'd2: value = 3'd7;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd4: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd6;
                5'd2: value = 3'd6;
                5'd3: value = 3'd6;
                5'd4: value = 3'd6;
                5'd5: value = 3'd6;
                5'd6: value = 3'd6;
                5'd7: value = 3'd6;
                5'd8: value = 3'd6;
                5'd9: value = 3'd6;
                5'd10: value = 3'd6;
                5'd11: value = 3'd6;
                5'd12: value = 3'd6;
                5'd13: value = 3'd6;
                5'd14: value = 3'd6;
                5'd15: value = 3'd6;
                5'd16: value = 3'd6;
                5'd17: value = 3'd6;
                5'd18: value = 3'd6;
                5'd19: value = 3'd6;
                5'd20: value = 3'd6;
                5'd21: value = 3'd6;
                5'd22: value = 3'd6;
                5'd23: value = 3'd6;
                5'd24: value = 3'd6;
                5'd25: value = 3'd6;
                5'd26: value = 3'd6;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd5: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd4;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd6: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd4;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd4;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd7: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd6;
                5'd4: value = 3'd6;
                5'd5: value = 3'd6;
                5'd6: value = 3'd6;
                5'd7: value = 3'd6;
                5'd8: value = 3'd6;
                5'd9: value = 3'd6;
                5'd10: value = 3'd6;
                5'd11: value = 3'd6;
                5'd12: value = 3'd6;
                5'd13: value = 3'd6;
                5'd14: value = 3'd6;
                5'd15: value = 3'd6;
                5'd16: value = 3'd6;
                5'd17: value = 3'd6;
                5'd18: value = 3'd6;
                5'd19: value = 3'd6;
                5'd20: value = 3'd6;
                5'd21: value = 3'd6;
                5'd22: value = 3'd6;
                5'd23: value = 3'd6;
                5'd24: value = 3'd6;
                5'd25: value = 3'd6;
                5'd26: value = 3'd6;
                5'd27: value = 3'd6;
                5'd28: value = 3'd6;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd8: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd5;
                5'd4: value = 3'd5;
                5'd5: value = 3'd5;
                5'd6: value = 3'd5;
                5'd7: value = 3'd5;
                5'd8: value = 3'd5;
                5'd9: value = 3'd5;
                5'd10: value = 3'd5;
                5'd11: value = 3'd5;
                5'd12: value = 3'd5;
                5'd13: value = 3'd5;
                5'd14: value = 3'd5;
                5'd15: value = 3'd5;
                5'd16: value = 3'd5;
                5'd17: value = 3'd5;
                5'd18: value = 3'd5;
                5'd19: value = 3'd5;
                5'd20: value = 3'd5;
                5'd21: value = 3'd5;
                5'd22: value = 3'd5;
                5'd23: value = 3'd5;
                5'd24: value = 3'd5;
                5'd25: value = 3'd5;
                5'd26: value = 3'd5;
                5'd27: value = 3'd5;
                5'd28: value = 3'd5;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd9: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd4;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd10: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd4;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd4;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd11: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd3;
                5'd2: value = 3'd3;
                5'd3: value = 3'd3;
                5'd4: value = 3'd3;
                5'd5: value = 3'd3;
                5'd6: value = 3'd3;
                5'd7: value = 3'd3;
                5'd8: value = 3'd3;
                5'd9: value = 3'd3;
                5'd10: value = 3'd3;
                5'd11: value = 3'd3;
                5'd12: value = 3'd3;
                5'd13: value = 3'd3;
                5'd14: value = 3'd3;
                5'd15: value = 3'd3;
                5'd16: value = 3'd3;
                5'd17: value = 3'd3;
                5'd18: value = 3'd3;
                5'd19: value = 3'd3;
                5'd20: value = 3'd3;
                5'd21: value = 3'd3;
                5'd22: value = 3'd3;
                5'd23: value = 3'd3;
                5'd24: value = 3'd3;
                5'd25: value = 3'd3;
                5'd26: value = 3'd3;
                5'd27: value = 3'd4;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd12: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd2;
                5'd2: value = 3'd2;
                5'd3: value = 3'd2;
                5'd4: value = 3'd2;
                5'd5: value = 3'd2;
                5'd6: value = 3'd2;
                5'd7: value = 3'd2;
                5'd8: value = 3'd2;
                5'd9: value = 3'd2;
                5'd10: value = 3'd2;
                5'd11: value = 3'd2;
                5'd12: value = 3'd2;
                5'd13: value = 3'd2;
                5'd14: value = 3'd2;
                5'd15: value = 3'd2;
                5'd16: value = 3'd2;
                5'd17: value = 3'd2;
                5'd18: value = 3'd2;
                5'd19: value = 3'd2;
                5'd20: value = 3'd2;
                5'd21: value = 3'd2;
                5'd22: value = 3'd2;
                5'd23: value = 3'd2;
                5'd24: value = 3'd2;
                5'd25: value = 3'd2;
                5'd26: value = 3'd2;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd13: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd4;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd4;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd14: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd4;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd4;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd15: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd1;
                5'd4: value = 3'd1;
                5'd5: value = 3'd1;
                5'd6: value = 3'd1;
                5'd7: value = 3'd1;
                5'd8: value = 3'd1;
                5'd9: value = 3'd1;
                5'd10: value = 3'd1;
                5'd11: value = 3'd1;
                5'd12: value = 3'd1;
                5'd13: value = 3'd1;
                5'd14: value = 3'd1;
                5'd15: value = 3'd1;
                5'd16: value = 3'd1;
                5'd17: value = 3'd1;
                5'd18: value = 3'd1;
                5'd19: value = 3'd1;
                5'd20: value = 3'd1;
                5'd21: value = 3'd1;
                5'd22: value = 3'd1;
                5'd23: value = 3'd1;
                5'd24: value = 3'd1;
                5'd25: value = 3'd1;
                5'd26: value = 3'd1;
                5'd27: value = 3'd1;
                5'd28: value = 3'd1;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd16: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd17: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd18: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd19: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd20: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd21: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd22: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd23: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd24: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd25: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd26: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd4;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd27: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd0;
                5'd26: value = 3'd0;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd28: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd29: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd4;
                5'd22: value = 3'd4;
                5'd23: value = 3'd4;
                5'd24: value = 3'd4;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd30: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd4;
                5'd22: value = 3'd4;
                5'd23: value = 3'd4;
                5'd24: value = 3'd4;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd31: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd4;
                5'd22: value = 3'd4;
                5'd23: value = 3'd4;
                5'd24: value = 3'd4;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd32: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd4;
                5'd22: value = 3'd4;
                5'd23: value = 3'd4;
                5'd24: value = 3'd4;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd33: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd34: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd35: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd36: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd37: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd4;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd38: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd0;
                5'd2: value = 3'd0;
                5'd3: value = 3'd0;
                5'd4: value = 3'd0;
                5'd5: value = 3'd0;
                5'd6: value = 3'd0;
                5'd7: value = 3'd0;
                5'd8: value = 3'd0;
                5'd9: value = 3'd0;
                5'd10: value = 3'd0;
                5'd11: value = 3'd0;
                5'd12: value = 3'd0;
                5'd13: value = 3'd0;
                5'd14: value = 3'd0;
                5'd15: value = 3'd0;
                5'd16: value = 3'd0;
                5'd17: value = 3'd0;
                5'd18: value = 3'd0;
                5'd19: value = 3'd0;
                5'd20: value = 3'd0;
                5'd21: value = 3'd0;
                5'd22: value = 3'd0;
                5'd23: value = 3'd0;
                5'd24: value = 3'd0;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd0;
                5'd28: value = 3'd0;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        6'd39: begin
            case (y)
                5'd0: value = 3'd7;
                5'd1: value = 3'd7;
                5'd2: value = 3'd7;
                5'd3: value = 3'd7;
                5'd4: value = 3'd7;
                5'd5: value = 3'd7;
                5'd6: value = 3'd7;
                5'd7: value = 3'd7;
                5'd8: value = 3'd7;
                5'd9: value = 3'd7;
                5'd10: value = 3'd7;
                5'd11: value = 3'd7;
                5'd12: value = 3'd7;
                5'd13: value = 3'd7;
                5'd14: value = 3'd7;
                5'd15: value = 3'd7;
                5'd16: value = 3'd7;
                5'd17: value = 3'd7;
                5'd18: value = 3'd7;
                5'd19: value = 3'd7;
                5'd20: value = 3'd7;
                5'd21: value = 3'd7;
                5'd22: value = 3'd7;
                5'd23: value = 3'd7;
                5'd24: value = 3'd7;
                5'd25: value = 3'd7;
                5'd26: value = 3'd7;
                5'd27: value = 3'd7;
                5'd28: value = 3'd7;
                5'd29: value = 3'd7;
                default: value = 3'd0;
            endcase
        end
        default: value = 3'd0;
    endcase
endmodule
