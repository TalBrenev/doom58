module grid(clock, reset, x, y, write, in, out);
    // Global clock and reset
    input clock;
    input reset;

    // Coordinates for the grid, write enable (read if off), grid value
    input [5:0] x;
    input [4:0] y;
    input write;
    input [2:0] in;

    // 3-bit output of what's contained in the grid address at xy
    output [2:0] out;
    reg [2:0] out;

    // 1200 3-bit Registers to store 40x30 grid squares of data
    reg [2:0] x0y0;
    reg [2:0] x0y1;
    reg [2:0] x0y2;
    reg [2:0] x0y3;
    reg [2:0] x0y4;
    reg [2:0] x0y5;
    reg [2:0] x0y6;
    reg [2:0] x0y7;
    reg [2:0] x0y8;
    reg [2:0] x0y9;
    reg [2:0] x0y10;
    reg [2:0] x0y11;
    reg [2:0] x0y12;
    reg [2:0] x0y13;
    reg [2:0] x0y14;
    reg [2:0] x0y15;
    reg [2:0] x0y16;
    reg [2:0] x0y17;
    reg [2:0] x0y18;
    reg [2:0] x0y19;
    reg [2:0] x0y20;
    reg [2:0] x0y21;
    reg [2:0] x0y22;
    reg [2:0] x0y23;
    reg [2:0] x0y24;
    reg [2:0] x0y25;
    reg [2:0] x0y26;
    reg [2:0] x0y27;
    reg [2:0] x0y28;
    reg [2:0] x0y29;
    reg [2:0] x1y0;
    reg [2:0] x1y1;
    reg [2:0] x1y2;
    reg [2:0] x1y3;
    reg [2:0] x1y4;
    reg [2:0] x1y5;
    reg [2:0] x1y6;
    reg [2:0] x1y7;
    reg [2:0] x1y8;
    reg [2:0] x1y9;
    reg [2:0] x1y10;
    reg [2:0] x1y11;
    reg [2:0] x1y12;
    reg [2:0] x1y13;
    reg [2:0] x1y14;
    reg [2:0] x1y15;
    reg [2:0] x1y16;
    reg [2:0] x1y17;
    reg [2:0] x1y18;
    reg [2:0] x1y19;
    reg [2:0] x1y20;
    reg [2:0] x1y21;
    reg [2:0] x1y22;
    reg [2:0] x1y23;
    reg [2:0] x1y24;
    reg [2:0] x1y25;
    reg [2:0] x1y26;
    reg [2:0] x1y27;
    reg [2:0] x1y28;
    reg [2:0] x1y29;
    reg [2:0] x2y0;
    reg [2:0] x2y1;
    reg [2:0] x2y2;
    reg [2:0] x2y3;
    reg [2:0] x2y4;
    reg [2:0] x2y5;
    reg [2:0] x2y6;
    reg [2:0] x2y7;
    reg [2:0] x2y8;
    reg [2:0] x2y9;
    reg [2:0] x2y10;
    reg [2:0] x2y11;
    reg [2:0] x2y12;
    reg [2:0] x2y13;
    reg [2:0] x2y14;
    reg [2:0] x2y15;
    reg [2:0] x2y16;
    reg [2:0] x2y17;
    reg [2:0] x2y18;
    reg [2:0] x2y19;
    reg [2:0] x2y20;
    reg [2:0] x2y21;
    reg [2:0] x2y22;
    reg [2:0] x2y23;
    reg [2:0] x2y24;
    reg [2:0] x2y25;
    reg [2:0] x2y26;
    reg [2:0] x2y27;
    reg [2:0] x2y28;
    reg [2:0] x2y29;
    reg [2:0] x3y0;
    reg [2:0] x3y1;
    reg [2:0] x3y2;
    reg [2:0] x3y3;
    reg [2:0] x3y4;
    reg [2:0] x3y5;
    reg [2:0] x3y6;
    reg [2:0] x3y7;
    reg [2:0] x3y8;
    reg [2:0] x3y9;
    reg [2:0] x3y10;
    reg [2:0] x3y11;
    reg [2:0] x3y12;
    reg [2:0] x3y13;
    reg [2:0] x3y14;
    reg [2:0] x3y15;
    reg [2:0] x3y16;
    reg [2:0] x3y17;
    reg [2:0] x3y18;
    reg [2:0] x3y19;
    reg [2:0] x3y20;
    reg [2:0] x3y21;
    reg [2:0] x3y22;
    reg [2:0] x3y23;
    reg [2:0] x3y24;
    reg [2:0] x3y25;
    reg [2:0] x3y26;
    reg [2:0] x3y27;
    reg [2:0] x3y28;
    reg [2:0] x3y29;
    reg [2:0] x4y0;
    reg [2:0] x4y1;
    reg [2:0] x4y2;
    reg [2:0] x4y3;
    reg [2:0] x4y4;
    reg [2:0] x4y5;
    reg [2:0] x4y6;
    reg [2:0] x4y7;
    reg [2:0] x4y8;
    reg [2:0] x4y9;
    reg [2:0] x4y10;
    reg [2:0] x4y11;
    reg [2:0] x4y12;
    reg [2:0] x4y13;
    reg [2:0] x4y14;
    reg [2:0] x4y15;
    reg [2:0] x4y16;
    reg [2:0] x4y17;
    reg [2:0] x4y18;
    reg [2:0] x4y19;
    reg [2:0] x4y20;
    reg [2:0] x4y21;
    reg [2:0] x4y22;
    reg [2:0] x4y23;
    reg [2:0] x4y24;
    reg [2:0] x4y25;
    reg [2:0] x4y26;
    reg [2:0] x4y27;
    reg [2:0] x4y28;
    reg [2:0] x4y29;
    reg [2:0] x5y0;
    reg [2:0] x5y1;
    reg [2:0] x5y2;
    reg [2:0] x5y3;
    reg [2:0] x5y4;
    reg [2:0] x5y5;
    reg [2:0] x5y6;
    reg [2:0] x5y7;
    reg [2:0] x5y8;
    reg [2:0] x5y9;
    reg [2:0] x5y10;
    reg [2:0] x5y11;
    reg [2:0] x5y12;
    reg [2:0] x5y13;
    reg [2:0] x5y14;
    reg [2:0] x5y15;
    reg [2:0] x5y16;
    reg [2:0] x5y17;
    reg [2:0] x5y18;
    reg [2:0] x5y19;
    reg [2:0] x5y20;
    reg [2:0] x5y21;
    reg [2:0] x5y22;
    reg [2:0] x5y23;
    reg [2:0] x5y24;
    reg [2:0] x5y25;
    reg [2:0] x5y26;
    reg [2:0] x5y27;
    reg [2:0] x5y28;
    reg [2:0] x5y29;
    reg [2:0] x6y0;
    reg [2:0] x6y1;
    reg [2:0] x6y2;
    reg [2:0] x6y3;
    reg [2:0] x6y4;
    reg [2:0] x6y5;
    reg [2:0] x6y6;
    reg [2:0] x6y7;
    reg [2:0] x6y8;
    reg [2:0] x6y9;
    reg [2:0] x6y10;
    reg [2:0] x6y11;
    reg [2:0] x6y12;
    reg [2:0] x6y13;
    reg [2:0] x6y14;
    reg [2:0] x6y15;
    reg [2:0] x6y16;
    reg [2:0] x6y17;
    reg [2:0] x6y18;
    reg [2:0] x6y19;
    reg [2:0] x6y20;
    reg [2:0] x6y21;
    reg [2:0] x6y22;
    reg [2:0] x6y23;
    reg [2:0] x6y24;
    reg [2:0] x6y25;
    reg [2:0] x6y26;
    reg [2:0] x6y27;
    reg [2:0] x6y28;
    reg [2:0] x6y29;
    reg [2:0] x7y0;
    reg [2:0] x7y1;
    reg [2:0] x7y2;
    reg [2:0] x7y3;
    reg [2:0] x7y4;
    reg [2:0] x7y5;
    reg [2:0] x7y6;
    reg [2:0] x7y7;
    reg [2:0] x7y8;
    reg [2:0] x7y9;
    reg [2:0] x7y10;
    reg [2:0] x7y11;
    reg [2:0] x7y12;
    reg [2:0] x7y13;
    reg [2:0] x7y14;
    reg [2:0] x7y15;
    reg [2:0] x7y16;
    reg [2:0] x7y17;
    reg [2:0] x7y18;
    reg [2:0] x7y19;
    reg [2:0] x7y20;
    reg [2:0] x7y21;
    reg [2:0] x7y22;
    reg [2:0] x7y23;
    reg [2:0] x7y24;
    reg [2:0] x7y25;
    reg [2:0] x7y26;
    reg [2:0] x7y27;
    reg [2:0] x7y28;
    reg [2:0] x7y29;
    reg [2:0] x8y0;
    reg [2:0] x8y1;
    reg [2:0] x8y2;
    reg [2:0] x8y3;
    reg [2:0] x8y4;
    reg [2:0] x8y5;
    reg [2:0] x8y6;
    reg [2:0] x8y7;
    reg [2:0] x8y8;
    reg [2:0] x8y9;
    reg [2:0] x8y10;
    reg [2:0] x8y11;
    reg [2:0] x8y12;
    reg [2:0] x8y13;
    reg [2:0] x8y14;
    reg [2:0] x8y15;
    reg [2:0] x8y16;
    reg [2:0] x8y17;
    reg [2:0] x8y18;
    reg [2:0] x8y19;
    reg [2:0] x8y20;
    reg [2:0] x8y21;
    reg [2:0] x8y22;
    reg [2:0] x8y23;
    reg [2:0] x8y24;
    reg [2:0] x8y25;
    reg [2:0] x8y26;
    reg [2:0] x8y27;
    reg [2:0] x8y28;
    reg [2:0] x8y29;
    reg [2:0] x9y0;
    reg [2:0] x9y1;
    reg [2:0] x9y2;
    reg [2:0] x9y3;
    reg [2:0] x9y4;
    reg [2:0] x9y5;
    reg [2:0] x9y6;
    reg [2:0] x9y7;
    reg [2:0] x9y8;
    reg [2:0] x9y9;
    reg [2:0] x9y10;
    reg [2:0] x9y11;
    reg [2:0] x9y12;
    reg [2:0] x9y13;
    reg [2:0] x9y14;
    reg [2:0] x9y15;
    reg [2:0] x9y16;
    reg [2:0] x9y17;
    reg [2:0] x9y18;
    reg [2:0] x9y19;
    reg [2:0] x9y20;
    reg [2:0] x9y21;
    reg [2:0] x9y22;
    reg [2:0] x9y23;
    reg [2:0] x9y24;
    reg [2:0] x9y25;
    reg [2:0] x9y26;
    reg [2:0] x9y27;
    reg [2:0] x9y28;
    reg [2:0] x9y29;
    reg [2:0] x10y0;
    reg [2:0] x10y1;
    reg [2:0] x10y2;
    reg [2:0] x10y3;
    reg [2:0] x10y4;
    reg [2:0] x10y5;
    reg [2:0] x10y6;
    reg [2:0] x10y7;
    reg [2:0] x10y8;
    reg [2:0] x10y9;
    reg [2:0] x10y10;
    reg [2:0] x10y11;
    reg [2:0] x10y12;
    reg [2:0] x10y13;
    reg [2:0] x10y14;
    reg [2:0] x10y15;
    reg [2:0] x10y16;
    reg [2:0] x10y17;
    reg [2:0] x10y18;
    reg [2:0] x10y19;
    reg [2:0] x10y20;
    reg [2:0] x10y21;
    reg [2:0] x10y22;
    reg [2:0] x10y23;
    reg [2:0] x10y24;
    reg [2:0] x10y25;
    reg [2:0] x10y26;
    reg [2:0] x10y27;
    reg [2:0] x10y28;
    reg [2:0] x10y29;
    reg [2:0] x11y0;
    reg [2:0] x11y1;
    reg [2:0] x11y2;
    reg [2:0] x11y3;
    reg [2:0] x11y4;
    reg [2:0] x11y5;
    reg [2:0] x11y6;
    reg [2:0] x11y7;
    reg [2:0] x11y8;
    reg [2:0] x11y9;
    reg [2:0] x11y10;
    reg [2:0] x11y11;
    reg [2:0] x11y12;
    reg [2:0] x11y13;
    reg [2:0] x11y14;
    reg [2:0] x11y15;
    reg [2:0] x11y16;
    reg [2:0] x11y17;
    reg [2:0] x11y18;
    reg [2:0] x11y19;
    reg [2:0] x11y20;
    reg [2:0] x11y21;
    reg [2:0] x11y22;
    reg [2:0] x11y23;
    reg [2:0] x11y24;
    reg [2:0] x11y25;
    reg [2:0] x11y26;
    reg [2:0] x11y27;
    reg [2:0] x11y28;
    reg [2:0] x11y29;
    reg [2:0] x12y0;
    reg [2:0] x12y1;
    reg [2:0] x12y2;
    reg [2:0] x12y3;
    reg [2:0] x12y4;
    reg [2:0] x12y5;
    reg [2:0] x12y6;
    reg [2:0] x12y7;
    reg [2:0] x12y8;
    reg [2:0] x12y9;
    reg [2:0] x12y10;
    reg [2:0] x12y11;
    reg [2:0] x12y12;
    reg [2:0] x12y13;
    reg [2:0] x12y14;
    reg [2:0] x12y15;
    reg [2:0] x12y16;
    reg [2:0] x12y17;
    reg [2:0] x12y18;
    reg [2:0] x12y19;
    reg [2:0] x12y20;
    reg [2:0] x12y21;
    reg [2:0] x12y22;
    reg [2:0] x12y23;
    reg [2:0] x12y24;
    reg [2:0] x12y25;
    reg [2:0] x12y26;
    reg [2:0] x12y27;
    reg [2:0] x12y28;
    reg [2:0] x12y29;
    reg [2:0] x13y0;
    reg [2:0] x13y1;
    reg [2:0] x13y2;
    reg [2:0] x13y3;
    reg [2:0] x13y4;
    reg [2:0] x13y5;
    reg [2:0] x13y6;
    reg [2:0] x13y7;
    reg [2:0] x13y8;
    reg [2:0] x13y9;
    reg [2:0] x13y10;
    reg [2:0] x13y11;
    reg [2:0] x13y12;
    reg [2:0] x13y13;
    reg [2:0] x13y14;
    reg [2:0] x13y15;
    reg [2:0] x13y16;
    reg [2:0] x13y17;
    reg [2:0] x13y18;
    reg [2:0] x13y19;
    reg [2:0] x13y20;
    reg [2:0] x13y21;
    reg [2:0] x13y22;
    reg [2:0] x13y23;
    reg [2:0] x13y24;
    reg [2:0] x13y25;
    reg [2:0] x13y26;
    reg [2:0] x13y27;
    reg [2:0] x13y28;
    reg [2:0] x13y29;
    reg [2:0] x14y0;
    reg [2:0] x14y1;
    reg [2:0] x14y2;
    reg [2:0] x14y3;
    reg [2:0] x14y4;
    reg [2:0] x14y5;
    reg [2:0] x14y6;
    reg [2:0] x14y7;
    reg [2:0] x14y8;
    reg [2:0] x14y9;
    reg [2:0] x14y10;
    reg [2:0] x14y11;
    reg [2:0] x14y12;
    reg [2:0] x14y13;
    reg [2:0] x14y14;
    reg [2:0] x14y15;
    reg [2:0] x14y16;
    reg [2:0] x14y17;
    reg [2:0] x14y18;
    reg [2:0] x14y19;
    reg [2:0] x14y20;
    reg [2:0] x14y21;
    reg [2:0] x14y22;
    reg [2:0] x14y23;
    reg [2:0] x14y24;
    reg [2:0] x14y25;
    reg [2:0] x14y26;
    reg [2:0] x14y27;
    reg [2:0] x14y28;
    reg [2:0] x14y29;
    reg [2:0] x15y0;
    reg [2:0] x15y1;
    reg [2:0] x15y2;
    reg [2:0] x15y3;
    reg [2:0] x15y4;
    reg [2:0] x15y5;
    reg [2:0] x15y6;
    reg [2:0] x15y7;
    reg [2:0] x15y8;
    reg [2:0] x15y9;
    reg [2:0] x15y10;
    reg [2:0] x15y11;
    reg [2:0] x15y12;
    reg [2:0] x15y13;
    reg [2:0] x15y14;
    reg [2:0] x15y15;
    reg [2:0] x15y16;
    reg [2:0] x15y17;
    reg [2:0] x15y18;
    reg [2:0] x15y19;
    reg [2:0] x15y20;
    reg [2:0] x15y21;
    reg [2:0] x15y22;
    reg [2:0] x15y23;
    reg [2:0] x15y24;
    reg [2:0] x15y25;
    reg [2:0] x15y26;
    reg [2:0] x15y27;
    reg [2:0] x15y28;
    reg [2:0] x15y29;
    reg [2:0] x16y0;
    reg [2:0] x16y1;
    reg [2:0] x16y2;
    reg [2:0] x16y3;
    reg [2:0] x16y4;
    reg [2:0] x16y5;
    reg [2:0] x16y6;
    reg [2:0] x16y7;
    reg [2:0] x16y8;
    reg [2:0] x16y9;
    reg [2:0] x16y10;
    reg [2:0] x16y11;
    reg [2:0] x16y12;
    reg [2:0] x16y13;
    reg [2:0] x16y14;
    reg [2:0] x16y15;
    reg [2:0] x16y16;
    reg [2:0] x16y17;
    reg [2:0] x16y18;
    reg [2:0] x16y19;
    reg [2:0] x16y20;
    reg [2:0] x16y21;
    reg [2:0] x16y22;
    reg [2:0] x16y23;
    reg [2:0] x16y24;
    reg [2:0] x16y25;
    reg [2:0] x16y26;
    reg [2:0] x16y27;
    reg [2:0] x16y28;
    reg [2:0] x16y29;
    reg [2:0] x17y0;
    reg [2:0] x17y1;
    reg [2:0] x17y2;
    reg [2:0] x17y3;
    reg [2:0] x17y4;
    reg [2:0] x17y5;
    reg [2:0] x17y6;
    reg [2:0] x17y7;
    reg [2:0] x17y8;
    reg [2:0] x17y9;
    reg [2:0] x17y10;
    reg [2:0] x17y11;
    reg [2:0] x17y12;
    reg [2:0] x17y13;
    reg [2:0] x17y14;
    reg [2:0] x17y15;
    reg [2:0] x17y16;
    reg [2:0] x17y17;
    reg [2:0] x17y18;
    reg [2:0] x17y19;
    reg [2:0] x17y20;
    reg [2:0] x17y21;
    reg [2:0] x17y22;
    reg [2:0] x17y23;
    reg [2:0] x17y24;
    reg [2:0] x17y25;
    reg [2:0] x17y26;
    reg [2:0] x17y27;
    reg [2:0] x17y28;
    reg [2:0] x17y29;
    reg [2:0] x18y0;
    reg [2:0] x18y1;
    reg [2:0] x18y2;
    reg [2:0] x18y3;
    reg [2:0] x18y4;
    reg [2:0] x18y5;
    reg [2:0] x18y6;
    reg [2:0] x18y7;
    reg [2:0] x18y8;
    reg [2:0] x18y9;
    reg [2:0] x18y10;
    reg [2:0] x18y11;
    reg [2:0] x18y12;
    reg [2:0] x18y13;
    reg [2:0] x18y14;
    reg [2:0] x18y15;
    reg [2:0] x18y16;
    reg [2:0] x18y17;
    reg [2:0] x18y18;
    reg [2:0] x18y19;
    reg [2:0] x18y20;
    reg [2:0] x18y21;
    reg [2:0] x18y22;
    reg [2:0] x18y23;
    reg [2:0] x18y24;
    reg [2:0] x18y25;
    reg [2:0] x18y26;
    reg [2:0] x18y27;
    reg [2:0] x18y28;
    reg [2:0] x18y29;
    reg [2:0] x19y0;
    reg [2:0] x19y1;
    reg [2:0] x19y2;
    reg [2:0] x19y3;
    reg [2:0] x19y4;
    reg [2:0] x19y5;
    reg [2:0] x19y6;
    reg [2:0] x19y7;
    reg [2:0] x19y8;
    reg [2:0] x19y9;
    reg [2:0] x19y10;
    reg [2:0] x19y11;
    reg [2:0] x19y12;
    reg [2:0] x19y13;
    reg [2:0] x19y14;
    reg [2:0] x19y15;
    reg [2:0] x19y16;
    reg [2:0] x19y17;
    reg [2:0] x19y18;
    reg [2:0] x19y19;
    reg [2:0] x19y20;
    reg [2:0] x19y21;
    reg [2:0] x19y22;
    reg [2:0] x19y23;
    reg [2:0] x19y24;
    reg [2:0] x19y25;
    reg [2:0] x19y26;
    reg [2:0] x19y27;
    reg [2:0] x19y28;
    reg [2:0] x19y29;
    reg [2:0] x20y0;
    reg [2:0] x20y1;
    reg [2:0] x20y2;
    reg [2:0] x20y3;
    reg [2:0] x20y4;
    reg [2:0] x20y5;
    reg [2:0] x20y6;
    reg [2:0] x20y7;
    reg [2:0] x20y8;
    reg [2:0] x20y9;
    reg [2:0] x20y10;
    reg [2:0] x20y11;
    reg [2:0] x20y12;
    reg [2:0] x20y13;
    reg [2:0] x20y14;
    reg [2:0] x20y15;
    reg [2:0] x20y16;
    reg [2:0] x20y17;
    reg [2:0] x20y18;
    reg [2:0] x20y19;
    reg [2:0] x20y20;
    reg [2:0] x20y21;
    reg [2:0] x20y22;
    reg [2:0] x20y23;
    reg [2:0] x20y24;
    reg [2:0] x20y25;
    reg [2:0] x20y26;
    reg [2:0] x20y27;
    reg [2:0] x20y28;
    reg [2:0] x20y29;
    reg [2:0] x21y0;
    reg [2:0] x21y1;
    reg [2:0] x21y2;
    reg [2:0] x21y3;
    reg [2:0] x21y4;
    reg [2:0] x21y5;
    reg [2:0] x21y6;
    reg [2:0] x21y7;
    reg [2:0] x21y8;
    reg [2:0] x21y9;
    reg [2:0] x21y10;
    reg [2:0] x21y11;
    reg [2:0] x21y12;
    reg [2:0] x21y13;
    reg [2:0] x21y14;
    reg [2:0] x21y15;
    reg [2:0] x21y16;
    reg [2:0] x21y17;
    reg [2:0] x21y18;
    reg [2:0] x21y19;
    reg [2:0] x21y20;
    reg [2:0] x21y21;
    reg [2:0] x21y22;
    reg [2:0] x21y23;
    reg [2:0] x21y24;
    reg [2:0] x21y25;
    reg [2:0] x21y26;
    reg [2:0] x21y27;
    reg [2:0] x21y28;
    reg [2:0] x21y29;
    reg [2:0] x22y0;
    reg [2:0] x22y1;
    reg [2:0] x22y2;
    reg [2:0] x22y3;
    reg [2:0] x22y4;
    reg [2:0] x22y5;
    reg [2:0] x22y6;
    reg [2:0] x22y7;
    reg [2:0] x22y8;
    reg [2:0] x22y9;
    reg [2:0] x22y10;
    reg [2:0] x22y11;
    reg [2:0] x22y12;
    reg [2:0] x22y13;
    reg [2:0] x22y14;
    reg [2:0] x22y15;
    reg [2:0] x22y16;
    reg [2:0] x22y17;
    reg [2:0] x22y18;
    reg [2:0] x22y19;
    reg [2:0] x22y20;
    reg [2:0] x22y21;
    reg [2:0] x22y22;
    reg [2:0] x22y23;
    reg [2:0] x22y24;
    reg [2:0] x22y25;
    reg [2:0] x22y26;
    reg [2:0] x22y27;
    reg [2:0] x22y28;
    reg [2:0] x22y29;
    reg [2:0] x23y0;
    reg [2:0] x23y1;
    reg [2:0] x23y2;
    reg [2:0] x23y3;
    reg [2:0] x23y4;
    reg [2:0] x23y5;
    reg [2:0] x23y6;
    reg [2:0] x23y7;
    reg [2:0] x23y8;
    reg [2:0] x23y9;
    reg [2:0] x23y10;
    reg [2:0] x23y11;
    reg [2:0] x23y12;
    reg [2:0] x23y13;
    reg [2:0] x23y14;
    reg [2:0] x23y15;
    reg [2:0] x23y16;
    reg [2:0] x23y17;
    reg [2:0] x23y18;
    reg [2:0] x23y19;
    reg [2:0] x23y20;
    reg [2:0] x23y21;
    reg [2:0] x23y22;
    reg [2:0] x23y23;
    reg [2:0] x23y24;
    reg [2:0] x23y25;
    reg [2:0] x23y26;
    reg [2:0] x23y27;
    reg [2:0] x23y28;
    reg [2:0] x23y29;
    reg [2:0] x24y0;
    reg [2:0] x24y1;
    reg [2:0] x24y2;
    reg [2:0] x24y3;
    reg [2:0] x24y4;
    reg [2:0] x24y5;
    reg [2:0] x24y6;
    reg [2:0] x24y7;
    reg [2:0] x24y8;
    reg [2:0] x24y9;
    reg [2:0] x24y10;
    reg [2:0] x24y11;
    reg [2:0] x24y12;
    reg [2:0] x24y13;
    reg [2:0] x24y14;
    reg [2:0] x24y15;
    reg [2:0] x24y16;
    reg [2:0] x24y17;
    reg [2:0] x24y18;
    reg [2:0] x24y19;
    reg [2:0] x24y20;
    reg [2:0] x24y21;
    reg [2:0] x24y22;
    reg [2:0] x24y23;
    reg [2:0] x24y24;
    reg [2:0] x24y25;
    reg [2:0] x24y26;
    reg [2:0] x24y27;
    reg [2:0] x24y28;
    reg [2:0] x24y29;
    reg [2:0] x25y0;
    reg [2:0] x25y1;
    reg [2:0] x25y2;
    reg [2:0] x25y3;
    reg [2:0] x25y4;
    reg [2:0] x25y5;
    reg [2:0] x25y6;
    reg [2:0] x25y7;
    reg [2:0] x25y8;
    reg [2:0] x25y9;
    reg [2:0] x25y10;
    reg [2:0] x25y11;
    reg [2:0] x25y12;
    reg [2:0] x25y13;
    reg [2:0] x25y14;
    reg [2:0] x25y15;
    reg [2:0] x25y16;
    reg [2:0] x25y17;
    reg [2:0] x25y18;
    reg [2:0] x25y19;
    reg [2:0] x25y20;
    reg [2:0] x25y21;
    reg [2:0] x25y22;
    reg [2:0] x25y23;
    reg [2:0] x25y24;
    reg [2:0] x25y25;
    reg [2:0] x25y26;
    reg [2:0] x25y27;
    reg [2:0] x25y28;
    reg [2:0] x25y29;
    reg [2:0] x26y0;
    reg [2:0] x26y1;
    reg [2:0] x26y2;
    reg [2:0] x26y3;
    reg [2:0] x26y4;
    reg [2:0] x26y5;
    reg [2:0] x26y6;
    reg [2:0] x26y7;
    reg [2:0] x26y8;
    reg [2:0] x26y9;
    reg [2:0] x26y10;
    reg [2:0] x26y11;
    reg [2:0] x26y12;
    reg [2:0] x26y13;
    reg [2:0] x26y14;
    reg [2:0] x26y15;
    reg [2:0] x26y16;
    reg [2:0] x26y17;
    reg [2:0] x26y18;
    reg [2:0] x26y19;
    reg [2:0] x26y20;
    reg [2:0] x26y21;
    reg [2:0] x26y22;
    reg [2:0] x26y23;
    reg [2:0] x26y24;
    reg [2:0] x26y25;
    reg [2:0] x26y26;
    reg [2:0] x26y27;
    reg [2:0] x26y28;
    reg [2:0] x26y29;
    reg [2:0] x27y0;
    reg [2:0] x27y1;
    reg [2:0] x27y2;
    reg [2:0] x27y3;
    reg [2:0] x27y4;
    reg [2:0] x27y5;
    reg [2:0] x27y6;
    reg [2:0] x27y7;
    reg [2:0] x27y8;
    reg [2:0] x27y9;
    reg [2:0] x27y10;
    reg [2:0] x27y11;
    reg [2:0] x27y12;
    reg [2:0] x27y13;
    reg [2:0] x27y14;
    reg [2:0] x27y15;
    reg [2:0] x27y16;
    reg [2:0] x27y17;
    reg [2:0] x27y18;
    reg [2:0] x27y19;
    reg [2:0] x27y20;
    reg [2:0] x27y21;
    reg [2:0] x27y22;
    reg [2:0] x27y23;
    reg [2:0] x27y24;
    reg [2:0] x27y25;
    reg [2:0] x27y26;
    reg [2:0] x27y27;
    reg [2:0] x27y28;
    reg [2:0] x27y29;
    reg [2:0] x28y0;
    reg [2:0] x28y1;
    reg [2:0] x28y2;
    reg [2:0] x28y3;
    reg [2:0] x28y4;
    reg [2:0] x28y5;
    reg [2:0] x28y6;
    reg [2:0] x28y7;
    reg [2:0] x28y8;
    reg [2:0] x28y9;
    reg [2:0] x28y10;
    reg [2:0] x28y11;
    reg [2:0] x28y12;
    reg [2:0] x28y13;
    reg [2:0] x28y14;
    reg [2:0] x28y15;
    reg [2:0] x28y16;
    reg [2:0] x28y17;
    reg [2:0] x28y18;
    reg [2:0] x28y19;
    reg [2:0] x28y20;
    reg [2:0] x28y21;
    reg [2:0] x28y22;
    reg [2:0] x28y23;
    reg [2:0] x28y24;
    reg [2:0] x28y25;
    reg [2:0] x28y26;
    reg [2:0] x28y27;
    reg [2:0] x28y28;
    reg [2:0] x28y29;
    reg [2:0] x29y0;
    reg [2:0] x29y1;
    reg [2:0] x29y2;
    reg [2:0] x29y3;
    reg [2:0] x29y4;
    reg [2:0] x29y5;
    reg [2:0] x29y6;
    reg [2:0] x29y7;
    reg [2:0] x29y8;
    reg [2:0] x29y9;
    reg [2:0] x29y10;
    reg [2:0] x29y11;
    reg [2:0] x29y12;
    reg [2:0] x29y13;
    reg [2:0] x29y14;
    reg [2:0] x29y15;
    reg [2:0] x29y16;
    reg [2:0] x29y17;
    reg [2:0] x29y18;
    reg [2:0] x29y19;
    reg [2:0] x29y20;
    reg [2:0] x29y21;
    reg [2:0] x29y22;
    reg [2:0] x29y23;
    reg [2:0] x29y24;
    reg [2:0] x29y25;
    reg [2:0] x29y26;
    reg [2:0] x29y27;
    reg [2:0] x29y28;
    reg [2:0] x29y29;
    reg [2:0] x30y0;
    reg [2:0] x30y1;
    reg [2:0] x30y2;
    reg [2:0] x30y3;
    reg [2:0] x30y4;
    reg [2:0] x30y5;
    reg [2:0] x30y6;
    reg [2:0] x30y7;
    reg [2:0] x30y8;
    reg [2:0] x30y9;
    reg [2:0] x30y10;
    reg [2:0] x30y11;
    reg [2:0] x30y12;
    reg [2:0] x30y13;
    reg [2:0] x30y14;
    reg [2:0] x30y15;
    reg [2:0] x30y16;
    reg [2:0] x30y17;
    reg [2:0] x30y18;
    reg [2:0] x30y19;
    reg [2:0] x30y20;
    reg [2:0] x30y21;
    reg [2:0] x30y22;
    reg [2:0] x30y23;
    reg [2:0] x30y24;
    reg [2:0] x30y25;
    reg [2:0] x30y26;
    reg [2:0] x30y27;
    reg [2:0] x30y28;
    reg [2:0] x30y29;
    reg [2:0] x31y0;
    reg [2:0] x31y1;
    reg [2:0] x31y2;
    reg [2:0] x31y3;
    reg [2:0] x31y4;
    reg [2:0] x31y5;
    reg [2:0] x31y6;
    reg [2:0] x31y7;
    reg [2:0] x31y8;
    reg [2:0] x31y9;
    reg [2:0] x31y10;
    reg [2:0] x31y11;
    reg [2:0] x31y12;
    reg [2:0] x31y13;
    reg [2:0] x31y14;
    reg [2:0] x31y15;
    reg [2:0] x31y16;
    reg [2:0] x31y17;
    reg [2:0] x31y18;
    reg [2:0] x31y19;
    reg [2:0] x31y20;
    reg [2:0] x31y21;
    reg [2:0] x31y22;
    reg [2:0] x31y23;
    reg [2:0] x31y24;
    reg [2:0] x31y25;
    reg [2:0] x31y26;
    reg [2:0] x31y27;
    reg [2:0] x31y28;
    reg [2:0] x31y29;
    reg [2:0] x32y0;
    reg [2:0] x32y1;
    reg [2:0] x32y2;
    reg [2:0] x32y3;
    reg [2:0] x32y4;
    reg [2:0] x32y5;
    reg [2:0] x32y6;
    reg [2:0] x32y7;
    reg [2:0] x32y8;
    reg [2:0] x32y9;
    reg [2:0] x32y10;
    reg [2:0] x32y11;
    reg [2:0] x32y12;
    reg [2:0] x32y13;
    reg [2:0] x32y14;
    reg [2:0] x32y15;
    reg [2:0] x32y16;
    reg [2:0] x32y17;
    reg [2:0] x32y18;
    reg [2:0] x32y19;
    reg [2:0] x32y20;
    reg [2:0] x32y21;
    reg [2:0] x32y22;
    reg [2:0] x32y23;
    reg [2:0] x32y24;
    reg [2:0] x32y25;
    reg [2:0] x32y26;
    reg [2:0] x32y27;
    reg [2:0] x32y28;
    reg [2:0] x32y29;
    reg [2:0] x33y0;
    reg [2:0] x33y1;
    reg [2:0] x33y2;
    reg [2:0] x33y3;
    reg [2:0] x33y4;
    reg [2:0] x33y5;
    reg [2:0] x33y6;
    reg [2:0] x33y7;
    reg [2:0] x33y8;
    reg [2:0] x33y9;
    reg [2:0] x33y10;
    reg [2:0] x33y11;
    reg [2:0] x33y12;
    reg [2:0] x33y13;
    reg [2:0] x33y14;
    reg [2:0] x33y15;
    reg [2:0] x33y16;
    reg [2:0] x33y17;
    reg [2:0] x33y18;
    reg [2:0] x33y19;
    reg [2:0] x33y20;
    reg [2:0] x33y21;
    reg [2:0] x33y22;
    reg [2:0] x33y23;
    reg [2:0] x33y24;
    reg [2:0] x33y25;
    reg [2:0] x33y26;
    reg [2:0] x33y27;
    reg [2:0] x33y28;
    reg [2:0] x33y29;
    reg [2:0] x34y0;
    reg [2:0] x34y1;
    reg [2:0] x34y2;
    reg [2:0] x34y3;
    reg [2:0] x34y4;
    reg [2:0] x34y5;
    reg [2:0] x34y6;
    reg [2:0] x34y7;
    reg [2:0] x34y8;
    reg [2:0] x34y9;
    reg [2:0] x34y10;
    reg [2:0] x34y11;
    reg [2:0] x34y12;
    reg [2:0] x34y13;
    reg [2:0] x34y14;
    reg [2:0] x34y15;
    reg [2:0] x34y16;
    reg [2:0] x34y17;
    reg [2:0] x34y18;
    reg [2:0] x34y19;
    reg [2:0] x34y20;
    reg [2:0] x34y21;
    reg [2:0] x34y22;
    reg [2:0] x34y23;
    reg [2:0] x34y24;
    reg [2:0] x34y25;
    reg [2:0] x34y26;
    reg [2:0] x34y27;
    reg [2:0] x34y28;
    reg [2:0] x34y29;
    reg [2:0] x35y0;
    reg [2:0] x35y1;
    reg [2:0] x35y2;
    reg [2:0] x35y3;
    reg [2:0] x35y4;
    reg [2:0] x35y5;
    reg [2:0] x35y6;
    reg [2:0] x35y7;
    reg [2:0] x35y8;
    reg [2:0] x35y9;
    reg [2:0] x35y10;
    reg [2:0] x35y11;
    reg [2:0] x35y12;
    reg [2:0] x35y13;
    reg [2:0] x35y14;
    reg [2:0] x35y15;
    reg [2:0] x35y16;
    reg [2:0] x35y17;
    reg [2:0] x35y18;
    reg [2:0] x35y19;
    reg [2:0] x35y20;
    reg [2:0] x35y21;
    reg [2:0] x35y22;
    reg [2:0] x35y23;
    reg [2:0] x35y24;
    reg [2:0] x35y25;
    reg [2:0] x35y26;
    reg [2:0] x35y27;
    reg [2:0] x35y28;
    reg [2:0] x35y29;
    reg [2:0] x36y0;
    reg [2:0] x36y1;
    reg [2:0] x36y2;
    reg [2:0] x36y3;
    reg [2:0] x36y4;
    reg [2:0] x36y5;
    reg [2:0] x36y6;
    reg [2:0] x36y7;
    reg [2:0] x36y8;
    reg [2:0] x36y9;
    reg [2:0] x36y10;
    reg [2:0] x36y11;
    reg [2:0] x36y12;
    reg [2:0] x36y13;
    reg [2:0] x36y14;
    reg [2:0] x36y15;
    reg [2:0] x36y16;
    reg [2:0] x36y17;
    reg [2:0] x36y18;
    reg [2:0] x36y19;
    reg [2:0] x36y20;
    reg [2:0] x36y21;
    reg [2:0] x36y22;
    reg [2:0] x36y23;
    reg [2:0] x36y24;
    reg [2:0] x36y25;
    reg [2:0] x36y26;
    reg [2:0] x36y27;
    reg [2:0] x36y28;
    reg [2:0] x36y29;
    reg [2:0] x37y0;
    reg [2:0] x37y1;
    reg [2:0] x37y2;
    reg [2:0] x37y3;
    reg [2:0] x37y4;
    reg [2:0] x37y5;
    reg [2:0] x37y6;
    reg [2:0] x37y7;
    reg [2:0] x37y8;
    reg [2:0] x37y9;
    reg [2:0] x37y10;
    reg [2:0] x37y11;
    reg [2:0] x37y12;
    reg [2:0] x37y13;
    reg [2:0] x37y14;
    reg [2:0] x37y15;
    reg [2:0] x37y16;
    reg [2:0] x37y17;
    reg [2:0] x37y18;
    reg [2:0] x37y19;
    reg [2:0] x37y20;
    reg [2:0] x37y21;
    reg [2:0] x37y22;
    reg [2:0] x37y23;
    reg [2:0] x37y24;
    reg [2:0] x37y25;
    reg [2:0] x37y26;
    reg [2:0] x37y27;
    reg [2:0] x37y28;
    reg [2:0] x37y29;
    reg [2:0] x38y0;
    reg [2:0] x38y1;
    reg [2:0] x38y2;
    reg [2:0] x38y3;
    reg [2:0] x38y4;
    reg [2:0] x38y5;
    reg [2:0] x38y6;
    reg [2:0] x38y7;
    reg [2:0] x38y8;
    reg [2:0] x38y9;
    reg [2:0] x38y10;
    reg [2:0] x38y11;
    reg [2:0] x38y12;
    reg [2:0] x38y13;
    reg [2:0] x38y14;
    reg [2:0] x38y15;
    reg [2:0] x38y16;
    reg [2:0] x38y17;
    reg [2:0] x38y18;
    reg [2:0] x38y19;
    reg [2:0] x38y20;
    reg [2:0] x38y21;
    reg [2:0] x38y22;
    reg [2:0] x38y23;
    reg [2:0] x38y24;
    reg [2:0] x38y25;
    reg [2:0] x38y26;
    reg [2:0] x38y27;
    reg [2:0] x38y28;
    reg [2:0] x38y29;
    reg [2:0] x39y0;
    reg [2:0] x39y1;
    reg [2:0] x39y2;
    reg [2:0] x39y3;
    reg [2:0] x39y4;
    reg [2:0] x39y5;
    reg [2:0] x39y6;
    reg [2:0] x39y7;
    reg [2:0] x39y8;
    reg [2:0] x39y9;
    reg [2:0] x39y10;
    reg [2:0] x39y11;
    reg [2:0] x39y12;
    reg [2:0] x39y13;
    reg [2:0] x39y14;
    reg [2:0] x39y15;
    reg [2:0] x39y16;
    reg [2:0] x39y17;
    reg [2:0] x39y18;
    reg [2:0] x39y19;
    reg [2:0] x39y20;
    reg [2:0] x39y21;
    reg [2:0] x39y22;
    reg [2:0] x39y23;
    reg [2:0] x39y24;
    reg [2:0] x39y25;
    reg [2:0] x39y26;
    reg [2:0] x39y27;
    reg [2:0] x39y28;
    reg [2:0] x39y29;

    // Assign 3-bit input to addresses when write enable on
    always @(posedge clock) begin
        if (write == 1) begin
            case (x)
                6'd0: begin
                    case (y)
                        5'd0: x0y0 = in;
                        5'd1: x0y1 = in;
                        5'd2: x0y2 = in;
                        5'd3: x0y3 = in;
                        5'd4: x0y4 = in;
                        5'd5: x0y5 = in;
                        5'd6: x0y6 = in;
                        5'd7: x0y7 = in;
                        5'd8: x0y8 = in;
                        5'd9: x0y9 = in;
                        5'd10: x0y10 = in;
                        5'd11: x0y11 = in;
                        5'd12: x0y12 = in;
                        5'd13: x0y13 = in;
                        5'd14: x0y14 = in;
                        5'd15: x0y15 = in;
                        5'd16: x0y16 = in;
                        5'd17: x0y17 = in;
                        5'd18: x0y18 = in;
                        5'd19: x0y19 = in;
                        5'd20: x0y20 = in;
                        5'd21: x0y21 = in;
                        5'd22: x0y22 = in;
                        5'd23: x0y23 = in;
                        5'd24: x0y24 = in;
                        5'd25: x0y25 = in;
                        5'd26: x0y26 = in;
                        5'd27: x0y27 = in;
                        5'd28: x0y28 = in;
                        5'd29: x0y29 = in;
                        default: ;
                    endcase
                end
                6'd1: begin
                    case (y)
                        5'd0: x1y0 = in;
                        5'd1: x1y1 = in;
                        5'd2: x1y2 = in;
                        5'd3: x1y3 = in;
                        5'd4: x1y4 = in;
                        5'd5: x1y5 = in;
                        5'd6: x1y6 = in;
                        5'd7: x1y7 = in;
                        5'd8: x1y8 = in;
                        5'd9: x1y9 = in;
                        5'd10: x1y10 = in;
                        5'd11: x1y11 = in;
                        5'd12: x1y12 = in;
                        5'd13: x1y13 = in;
                        5'd14: x1y14 = in;
                        5'd15: x1y15 = in;
                        5'd16: x1y16 = in;
                        5'd17: x1y17 = in;
                        5'd18: x1y18 = in;
                        5'd19: x1y19 = in;
                        5'd20: x1y20 = in;
                        5'd21: x1y21 = in;
                        5'd22: x1y22 = in;
                        5'd23: x1y23 = in;
                        5'd24: x1y24 = in;
                        5'd25: x1y25 = in;
                        5'd26: x1y26 = in;
                        5'd27: x1y27 = in;
                        5'd28: x1y28 = in;
                        5'd29: x1y29 = in;
                        default: ;
                    endcase
                end
                6'd2: begin
                    case (y)
                        5'd0: x2y0 = in;
                        5'd1: x2y1 = in;
                        5'd2: x2y2 = in;
                        5'd3: x2y3 = in;
                        5'd4: x2y4 = in;
                        5'd5: x2y5 = in;
                        5'd6: x2y6 = in;
                        5'd7: x2y7 = in;
                        5'd8: x2y8 = in;
                        5'd9: x2y9 = in;
                        5'd10: x2y10 = in;
                        5'd11: x2y11 = in;
                        5'd12: x2y12 = in;
                        5'd13: x2y13 = in;
                        5'd14: x2y14 = in;
                        5'd15: x2y15 = in;
                        5'd16: x2y16 = in;
                        5'd17: x2y17 = in;
                        5'd18: x2y18 = in;
                        5'd19: x2y19 = in;
                        5'd20: x2y20 = in;
                        5'd21: x2y21 = in;
                        5'd22: x2y22 = in;
                        5'd23: x2y23 = in;
                        5'd24: x2y24 = in;
                        5'd25: x2y25 = in;
                        5'd26: x2y26 = in;
                        5'd27: x2y27 = in;
                        5'd28: x2y28 = in;
                        5'd29: x2y29 = in;
                        default: ;
                    endcase
                end
                6'd3: begin
                    case (y)
                        5'd0: x3y0 = in;
                        5'd1: x3y1 = in;
                        5'd2: x3y2 = in;
                        5'd3: x3y3 = in;
                        5'd4: x3y4 = in;
                        5'd5: x3y5 = in;
                        5'd6: x3y6 = in;
                        5'd7: x3y7 = in;
                        5'd8: x3y8 = in;
                        5'd9: x3y9 = in;
                        5'd10: x3y10 = in;
                        5'd11: x3y11 = in;
                        5'd12: x3y12 = in;
                        5'd13: x3y13 = in;
                        5'd14: x3y14 = in;
                        5'd15: x3y15 = in;
                        5'd16: x3y16 = in;
                        5'd17: x3y17 = in;
                        5'd18: x3y18 = in;
                        5'd19: x3y19 = in;
                        5'd20: x3y20 = in;
                        5'd21: x3y21 = in;
                        5'd22: x3y22 = in;
                        5'd23: x3y23 = in;
                        5'd24: x3y24 = in;
                        5'd25: x3y25 = in;
                        5'd26: x3y26 = in;
                        5'd27: x3y27 = in;
                        5'd28: x3y28 = in;
                        5'd29: x3y29 = in;
                        default: ;
                    endcase
                end
                6'd4: begin
                    case (y)
                        5'd0: x4y0 = in;
                        5'd1: x4y1 = in;
                        5'd2: x4y2 = in;
                        5'd3: x4y3 = in;
                        5'd4: x4y4 = in;
                        5'd5: x4y5 = in;
                        5'd6: x4y6 = in;
                        5'd7: x4y7 = in;
                        5'd8: x4y8 = in;
                        5'd9: x4y9 = in;
                        5'd10: x4y10 = in;
                        5'd11: x4y11 = in;
                        5'd12: x4y12 = in;
                        5'd13: x4y13 = in;
                        5'd14: x4y14 = in;
                        5'd15: x4y15 = in;
                        5'd16: x4y16 = in;
                        5'd17: x4y17 = in;
                        5'd18: x4y18 = in;
                        5'd19: x4y19 = in;
                        5'd20: x4y20 = in;
                        5'd21: x4y21 = in;
                        5'd22: x4y22 = in;
                        5'd23: x4y23 = in;
                        5'd24: x4y24 = in;
                        5'd25: x4y25 = in;
                        5'd26: x4y26 = in;
                        5'd27: x4y27 = in;
                        5'd28: x4y28 = in;
                        5'd29: x4y29 = in;
                        default: ;
                    endcase
                end
                6'd5: begin
                    case (y)
                        5'd0: x5y0 = in;
                        5'd1: x5y1 = in;
                        5'd2: x5y2 = in;
                        5'd3: x5y3 = in;
                        5'd4: x5y4 = in;
                        5'd5: x5y5 = in;
                        5'd6: x5y6 = in;
                        5'd7: x5y7 = in;
                        5'd8: x5y8 = in;
                        5'd9: x5y9 = in;
                        5'd10: x5y10 = in;
                        5'd11: x5y11 = in;
                        5'd12: x5y12 = in;
                        5'd13: x5y13 = in;
                        5'd14: x5y14 = in;
                        5'd15: x5y15 = in;
                        5'd16: x5y16 = in;
                        5'd17: x5y17 = in;
                        5'd18: x5y18 = in;
                        5'd19: x5y19 = in;
                        5'd20: x5y20 = in;
                        5'd21: x5y21 = in;
                        5'd22: x5y22 = in;
                        5'd23: x5y23 = in;
                        5'd24: x5y24 = in;
                        5'd25: x5y25 = in;
                        5'd26: x5y26 = in;
                        5'd27: x5y27 = in;
                        5'd28: x5y28 = in;
                        5'd29: x5y29 = in;
                        default: ;
                    endcase
                end
                6'd6: begin
                    case (y)
                        5'd0: x6y0 = in;
                        5'd1: x6y1 = in;
                        5'd2: x6y2 = in;
                        5'd3: x6y3 = in;
                        5'd4: x6y4 = in;
                        5'd5: x6y5 = in;
                        5'd6: x6y6 = in;
                        5'd7: x6y7 = in;
                        5'd8: x6y8 = in;
                        5'd9: x6y9 = in;
                        5'd10: x6y10 = in;
                        5'd11: x6y11 = in;
                        5'd12: x6y12 = in;
                        5'd13: x6y13 = in;
                        5'd14: x6y14 = in;
                        5'd15: x6y15 = in;
                        5'd16: x6y16 = in;
                        5'd17: x6y17 = in;
                        5'd18: x6y18 = in;
                        5'd19: x6y19 = in;
                        5'd20: x6y20 = in;
                        5'd21: x6y21 = in;
                        5'd22: x6y22 = in;
                        5'd23: x6y23 = in;
                        5'd24: x6y24 = in;
                        5'd25: x6y25 = in;
                        5'd26: x6y26 = in;
                        5'd27: x6y27 = in;
                        5'd28: x6y28 = in;
                        5'd29: x6y29 = in;
                        default: ;
                    endcase
                end
                6'd7: begin
                    case (y)
                        5'd0: x7y0 = in;
                        5'd1: x7y1 = in;
                        5'd2: x7y2 = in;
                        5'd3: x7y3 = in;
                        5'd4: x7y4 = in;
                        5'd5: x7y5 = in;
                        5'd6: x7y6 = in;
                        5'd7: x7y7 = in;
                        5'd8: x7y8 = in;
                        5'd9: x7y9 = in;
                        5'd10: x7y10 = in;
                        5'd11: x7y11 = in;
                        5'd12: x7y12 = in;
                        5'd13: x7y13 = in;
                        5'd14: x7y14 = in;
                        5'd15: x7y15 = in;
                        5'd16: x7y16 = in;
                        5'd17: x7y17 = in;
                        5'd18: x7y18 = in;
                        5'd19: x7y19 = in;
                        5'd20: x7y20 = in;
                        5'd21: x7y21 = in;
                        5'd22: x7y22 = in;
                        5'd23: x7y23 = in;
                        5'd24: x7y24 = in;
                        5'd25: x7y25 = in;
                        5'd26: x7y26 = in;
                        5'd27: x7y27 = in;
                        5'd28: x7y28 = in;
                        5'd29: x7y29 = in;
                        default: ;
                    endcase
                end
                6'd8: begin
                    case (y)
                        5'd0: x8y0 = in;
                        5'd1: x8y1 = in;
                        5'd2: x8y2 = in;
                        5'd3: x8y3 = in;
                        5'd4: x8y4 = in;
                        5'd5: x8y5 = in;
                        5'd6: x8y6 = in;
                        5'd7: x8y7 = in;
                        5'd8: x8y8 = in;
                        5'd9: x8y9 = in;
                        5'd10: x8y10 = in;
                        5'd11: x8y11 = in;
                        5'd12: x8y12 = in;
                        5'd13: x8y13 = in;
                        5'd14: x8y14 = in;
                        5'd15: x8y15 = in;
                        5'd16: x8y16 = in;
                        5'd17: x8y17 = in;
                        5'd18: x8y18 = in;
                        5'd19: x8y19 = in;
                        5'd20: x8y20 = in;
                        5'd21: x8y21 = in;
                        5'd22: x8y22 = in;
                        5'd23: x8y23 = in;
                        5'd24: x8y24 = in;
                        5'd25: x8y25 = in;
                        5'd26: x8y26 = in;
                        5'd27: x8y27 = in;
                        5'd28: x8y28 = in;
                        5'd29: x8y29 = in;
                        default: ;
                    endcase
                end
                6'd9: begin
                    case (y)
                        5'd0: x9y0 = in;
                        5'd1: x9y1 = in;
                        5'd2: x9y2 = in;
                        5'd3: x9y3 = in;
                        5'd4: x9y4 = in;
                        5'd5: x9y5 = in;
                        5'd6: x9y6 = in;
                        5'd7: x9y7 = in;
                        5'd8: x9y8 = in;
                        5'd9: x9y9 = in;
                        5'd10: x9y10 = in;
                        5'd11: x9y11 = in;
                        5'd12: x9y12 = in;
                        5'd13: x9y13 = in;
                        5'd14: x9y14 = in;
                        5'd15: x9y15 = in;
                        5'd16: x9y16 = in;
                        5'd17: x9y17 = in;
                        5'd18: x9y18 = in;
                        5'd19: x9y19 = in;
                        5'd20: x9y20 = in;
                        5'd21: x9y21 = in;
                        5'd22: x9y22 = in;
                        5'd23: x9y23 = in;
                        5'd24: x9y24 = in;
                        5'd25: x9y25 = in;
                        5'd26: x9y26 = in;
                        5'd27: x9y27 = in;
                        5'd28: x9y28 = in;
                        5'd29: x9y29 = in;
                        default: ;
                    endcase
                end
                6'd10: begin
                    case (y)
                        5'd0: x10y0 = in;
                        5'd1: x10y1 = in;
                        5'd2: x10y2 = in;
                        5'd3: x10y3 = in;
                        5'd4: x10y4 = in;
                        5'd5: x10y5 = in;
                        5'd6: x10y6 = in;
                        5'd7: x10y7 = in;
                        5'd8: x10y8 = in;
                        5'd9: x10y9 = in;
                        5'd10: x10y10 = in;
                        5'd11: x10y11 = in;
                        5'd12: x10y12 = in;
                        5'd13: x10y13 = in;
                        5'd14: x10y14 = in;
                        5'd15: x10y15 = in;
                        5'd16: x10y16 = in;
                        5'd17: x10y17 = in;
                        5'd18: x10y18 = in;
                        5'd19: x10y19 = in;
                        5'd20: x10y20 = in;
                        5'd21: x10y21 = in;
                        5'd22: x10y22 = in;
                        5'd23: x10y23 = in;
                        5'd24: x10y24 = in;
                        5'd25: x10y25 = in;
                        5'd26: x10y26 = in;
                        5'd27: x10y27 = in;
                        5'd28: x10y28 = in;
                        5'd29: x10y29 = in;
                        default: ;
                    endcase
                end
                6'd11: begin
                    case (y)
                        5'd0: x11y0 = in;
                        5'd1: x11y1 = in;
                        5'd2: x11y2 = in;
                        5'd3: x11y3 = in;
                        5'd4: x11y4 = in;
                        5'd5: x11y5 = in;
                        5'd6: x11y6 = in;
                        5'd7: x11y7 = in;
                        5'd8: x11y8 = in;
                        5'd9: x11y9 = in;
                        5'd10: x11y10 = in;
                        5'd11: x11y11 = in;
                        5'd12: x11y12 = in;
                        5'd13: x11y13 = in;
                        5'd14: x11y14 = in;
                        5'd15: x11y15 = in;
                        5'd16: x11y16 = in;
                        5'd17: x11y17 = in;
                        5'd18: x11y18 = in;
                        5'd19: x11y19 = in;
                        5'd20: x11y20 = in;
                        5'd21: x11y21 = in;
                        5'd22: x11y22 = in;
                        5'd23: x11y23 = in;
                        5'd24: x11y24 = in;
                        5'd25: x11y25 = in;
                        5'd26: x11y26 = in;
                        5'd27: x11y27 = in;
                        5'd28: x11y28 = in;
                        5'd29: x11y29 = in;
                        default: ;
                    endcase
                end
                6'd12: begin
                    case (y)
                        5'd0: x12y0 = in;
                        5'd1: x12y1 = in;
                        5'd2: x12y2 = in;
                        5'd3: x12y3 = in;
                        5'd4: x12y4 = in;
                        5'd5: x12y5 = in;
                        5'd6: x12y6 = in;
                        5'd7: x12y7 = in;
                        5'd8: x12y8 = in;
                        5'd9: x12y9 = in;
                        5'd10: x12y10 = in;
                        5'd11: x12y11 = in;
                        5'd12: x12y12 = in;
                        5'd13: x12y13 = in;
                        5'd14: x12y14 = in;
                        5'd15: x12y15 = in;
                        5'd16: x12y16 = in;
                        5'd17: x12y17 = in;
                        5'd18: x12y18 = in;
                        5'd19: x12y19 = in;
                        5'd20: x12y20 = in;
                        5'd21: x12y21 = in;
                        5'd22: x12y22 = in;
                        5'd23: x12y23 = in;
                        5'd24: x12y24 = in;
                        5'd25: x12y25 = in;
                        5'd26: x12y26 = in;
                        5'd27: x12y27 = in;
                        5'd28: x12y28 = in;
                        5'd29: x12y29 = in;
                        default: ;
                    endcase
                end
                6'd13: begin
                    case (y)
                        5'd0: x13y0 = in;
                        5'd1: x13y1 = in;
                        5'd2: x13y2 = in;
                        5'd3: x13y3 = in;
                        5'd4: x13y4 = in;
                        5'd5: x13y5 = in;
                        5'd6: x13y6 = in;
                        5'd7: x13y7 = in;
                        5'd8: x13y8 = in;
                        5'd9: x13y9 = in;
                        5'd10: x13y10 = in;
                        5'd11: x13y11 = in;
                        5'd12: x13y12 = in;
                        5'd13: x13y13 = in;
                        5'd14: x13y14 = in;
                        5'd15: x13y15 = in;
                        5'd16: x13y16 = in;
                        5'd17: x13y17 = in;
                        5'd18: x13y18 = in;
                        5'd19: x13y19 = in;
                        5'd20: x13y20 = in;
                        5'd21: x13y21 = in;
                        5'd22: x13y22 = in;
                        5'd23: x13y23 = in;
                        5'd24: x13y24 = in;
                        5'd25: x13y25 = in;
                        5'd26: x13y26 = in;
                        5'd27: x13y27 = in;
                        5'd28: x13y28 = in;
                        5'd29: x13y29 = in;
                        default: ;
                    endcase
                end
                6'd14: begin
                    case (y)
                        5'd0: x14y0 = in;
                        5'd1: x14y1 = in;
                        5'd2: x14y2 = in;
                        5'd3: x14y3 = in;
                        5'd4: x14y4 = in;
                        5'd5: x14y5 = in;
                        5'd6: x14y6 = in;
                        5'd7: x14y7 = in;
                        5'd8: x14y8 = in;
                        5'd9: x14y9 = in;
                        5'd10: x14y10 = in;
                        5'd11: x14y11 = in;
                        5'd12: x14y12 = in;
                        5'd13: x14y13 = in;
                        5'd14: x14y14 = in;
                        5'd15: x14y15 = in;
                        5'd16: x14y16 = in;
                        5'd17: x14y17 = in;
                        5'd18: x14y18 = in;
                        5'd19: x14y19 = in;
                        5'd20: x14y20 = in;
                        5'd21: x14y21 = in;
                        5'd22: x14y22 = in;
                        5'd23: x14y23 = in;
                        5'd24: x14y24 = in;
                        5'd25: x14y25 = in;
                        5'd26: x14y26 = in;
                        5'd27: x14y27 = in;
                        5'd28: x14y28 = in;
                        5'd29: x14y29 = in;
                        default: ;
                    endcase
                end
                6'd15: begin
                    case (y)
                        5'd0: x15y0 = in;
                        5'd1: x15y1 = in;
                        5'd2: x15y2 = in;
                        5'd3: x15y3 = in;
                        5'd4: x15y4 = in;
                        5'd5: x15y5 = in;
                        5'd6: x15y6 = in;
                        5'd7: x15y7 = in;
                        5'd8: x15y8 = in;
                        5'd9: x15y9 = in;
                        5'd10: x15y10 = in;
                        5'd11: x15y11 = in;
                        5'd12: x15y12 = in;
                        5'd13: x15y13 = in;
                        5'd14: x15y14 = in;
                        5'd15: x15y15 = in;
                        5'd16: x15y16 = in;
                        5'd17: x15y17 = in;
                        5'd18: x15y18 = in;
                        5'd19: x15y19 = in;
                        5'd20: x15y20 = in;
                        5'd21: x15y21 = in;
                        5'd22: x15y22 = in;
                        5'd23: x15y23 = in;
                        5'd24: x15y24 = in;
                        5'd25: x15y25 = in;
                        5'd26: x15y26 = in;
                        5'd27: x15y27 = in;
                        5'd28: x15y28 = in;
                        5'd29: x15y29 = in;
                        default: ;
                    endcase
                end
                6'd16: begin
                    case (y)
                        5'd0: x16y0 = in;
                        5'd1: x16y1 = in;
                        5'd2: x16y2 = in;
                        5'd3: x16y3 = in;
                        5'd4: x16y4 = in;
                        5'd5: x16y5 = in;
                        5'd6: x16y6 = in;
                        5'd7: x16y7 = in;
                        5'd8: x16y8 = in;
                        5'd9: x16y9 = in;
                        5'd10: x16y10 = in;
                        5'd11: x16y11 = in;
                        5'd12: x16y12 = in;
                        5'd13: x16y13 = in;
                        5'd14: x16y14 = in;
                        5'd15: x16y15 = in;
                        5'd16: x16y16 = in;
                        5'd17: x16y17 = in;
                        5'd18: x16y18 = in;
                        5'd19: x16y19 = in;
                        5'd20: x16y20 = in;
                        5'd21: x16y21 = in;
                        5'd22: x16y22 = in;
                        5'd23: x16y23 = in;
                        5'd24: x16y24 = in;
                        5'd25: x16y25 = in;
                        5'd26: x16y26 = in;
                        5'd27: x16y27 = in;
                        5'd28: x16y28 = in;
                        5'd29: x16y29 = in;
                        default: ;
                    endcase
                end
                6'd17: begin
                    case (y)
                        5'd0: x17y0 = in;
                        5'd1: x17y1 = in;
                        5'd2: x17y2 = in;
                        5'd3: x17y3 = in;
                        5'd4: x17y4 = in;
                        5'd5: x17y5 = in;
                        5'd6: x17y6 = in;
                        5'd7: x17y7 = in;
                        5'd8: x17y8 = in;
                        5'd9: x17y9 = in;
                        5'd10: x17y10 = in;
                        5'd11: x17y11 = in;
                        5'd12: x17y12 = in;
                        5'd13: x17y13 = in;
                        5'd14: x17y14 = in;
                        5'd15: x17y15 = in;
                        5'd16: x17y16 = in;
                        5'd17: x17y17 = in;
                        5'd18: x17y18 = in;
                        5'd19: x17y19 = in;
                        5'd20: x17y20 = in;
                        5'd21: x17y21 = in;
                        5'd22: x17y22 = in;
                        5'd23: x17y23 = in;
                        5'd24: x17y24 = in;
                        5'd25: x17y25 = in;
                        5'd26: x17y26 = in;
                        5'd27: x17y27 = in;
                        5'd28: x17y28 = in;
                        5'd29: x17y29 = in;
                        default: ;
                    endcase
                end
                6'd18: begin
                    case (y)
                        5'd0: x18y0 = in;
                        5'd1: x18y1 = in;
                        5'd2: x18y2 = in;
                        5'd3: x18y3 = in;
                        5'd4: x18y4 = in;
                        5'd5: x18y5 = in;
                        5'd6: x18y6 = in;
                        5'd7: x18y7 = in;
                        5'd8: x18y8 = in;
                        5'd9: x18y9 = in;
                        5'd10: x18y10 = in;
                        5'd11: x18y11 = in;
                        5'd12: x18y12 = in;
                        5'd13: x18y13 = in;
                        5'd14: x18y14 = in;
                        5'd15: x18y15 = in;
                        5'd16: x18y16 = in;
                        5'd17: x18y17 = in;
                        5'd18: x18y18 = in;
                        5'd19: x18y19 = in;
                        5'd20: x18y20 = in;
                        5'd21: x18y21 = in;
                        5'd22: x18y22 = in;
                        5'd23: x18y23 = in;
                        5'd24: x18y24 = in;
                        5'd25: x18y25 = in;
                        5'd26: x18y26 = in;
                        5'd27: x18y27 = in;
                        5'd28: x18y28 = in;
                        5'd29: x18y29 = in;
                        default: ;
                    endcase
                end
                6'd19: begin
                    case (y)
                        5'd0: x19y0 = in;
                        5'd1: x19y1 = in;
                        5'd2: x19y2 = in;
                        5'd3: x19y3 = in;
                        5'd4: x19y4 = in;
                        5'd5: x19y5 = in;
                        5'd6: x19y6 = in;
                        5'd7: x19y7 = in;
                        5'd8: x19y8 = in;
                        5'd9: x19y9 = in;
                        5'd10: x19y10 = in;
                        5'd11: x19y11 = in;
                        5'd12: x19y12 = in;
                        5'd13: x19y13 = in;
                        5'd14: x19y14 = in;
                        5'd15: x19y15 = in;
                        5'd16: x19y16 = in;
                        5'd17: x19y17 = in;
                        5'd18: x19y18 = in;
                        5'd19: x19y19 = in;
                        5'd20: x19y20 = in;
                        5'd21: x19y21 = in;
                        5'd22: x19y22 = in;
                        5'd23: x19y23 = in;
                        5'd24: x19y24 = in;
                        5'd25: x19y25 = in;
                        5'd26: x19y26 = in;
                        5'd27: x19y27 = in;
                        5'd28: x19y28 = in;
                        5'd29: x19y29 = in;
                        default: ;
                    endcase
                end
                6'd20: begin
                    case (y)
                        5'd0: x20y0 = in;
                        5'd1: x20y1 = in;
                        5'd2: x20y2 = in;
                        5'd3: x20y3 = in;
                        5'd4: x20y4 = in;
                        5'd5: x20y5 = in;
                        5'd6: x20y6 = in;
                        5'd7: x20y7 = in;
                        5'd8: x20y8 = in;
                        5'd9: x20y9 = in;
                        5'd10: x20y10 = in;
                        5'd11: x20y11 = in;
                        5'd12: x20y12 = in;
                        5'd13: x20y13 = in;
                        5'd14: x20y14 = in;
                        5'd15: x20y15 = in;
                        5'd16: x20y16 = in;
                        5'd17: x20y17 = in;
                        5'd18: x20y18 = in;
                        5'd19: x20y19 = in;
                        5'd20: x20y20 = in;
                        5'd21: x20y21 = in;
                        5'd22: x20y22 = in;
                        5'd23: x20y23 = in;
                        5'd24: x20y24 = in;
                        5'd25: x20y25 = in;
                        5'd26: x20y26 = in;
                        5'd27: x20y27 = in;
                        5'd28: x20y28 = in;
                        5'd29: x20y29 = in;
                        default: ;
                    endcase
                end
                6'd21: begin
                    case (y)
                        5'd0: x21y0 = in;
                        5'd1: x21y1 = in;
                        5'd2: x21y2 = in;
                        5'd3: x21y3 = in;
                        5'd4: x21y4 = in;
                        5'd5: x21y5 = in;
                        5'd6: x21y6 = in;
                        5'd7: x21y7 = in;
                        5'd8: x21y8 = in;
                        5'd9: x21y9 = in;
                        5'd10: x21y10 = in;
                        5'd11: x21y11 = in;
                        5'd12: x21y12 = in;
                        5'd13: x21y13 = in;
                        5'd14: x21y14 = in;
                        5'd15: x21y15 = in;
                        5'd16: x21y16 = in;
                        5'd17: x21y17 = in;
                        5'd18: x21y18 = in;
                        5'd19: x21y19 = in;
                        5'd20: x21y20 = in;
                        5'd21: x21y21 = in;
                        5'd22: x21y22 = in;
                        5'd23: x21y23 = in;
                        5'd24: x21y24 = in;
                        5'd25: x21y25 = in;
                        5'd26: x21y26 = in;
                        5'd27: x21y27 = in;
                        5'd28: x21y28 = in;
                        5'd29: x21y29 = in;
                        default: ;
                    endcase
                end
                6'd22: begin
                    case (y)
                        5'd0: x22y0 = in;
                        5'd1: x22y1 = in;
                        5'd2: x22y2 = in;
                        5'd3: x22y3 = in;
                        5'd4: x22y4 = in;
                        5'd5: x22y5 = in;
                        5'd6: x22y6 = in;
                        5'd7: x22y7 = in;
                        5'd8: x22y8 = in;
                        5'd9: x22y9 = in;
                        5'd10: x22y10 = in;
                        5'd11: x22y11 = in;
                        5'd12: x22y12 = in;
                        5'd13: x22y13 = in;
                        5'd14: x22y14 = in;
                        5'd15: x22y15 = in;
                        5'd16: x22y16 = in;
                        5'd17: x22y17 = in;
                        5'd18: x22y18 = in;
                        5'd19: x22y19 = in;
                        5'd20: x22y20 = in;
                        5'd21: x22y21 = in;
                        5'd22: x22y22 = in;
                        5'd23: x22y23 = in;
                        5'd24: x22y24 = in;
                        5'd25: x22y25 = in;
                        5'd26: x22y26 = in;
                        5'd27: x22y27 = in;
                        5'd28: x22y28 = in;
                        5'd29: x22y29 = in;
                        default: ;
                    endcase
                end
                6'd23: begin
                    case (y)
                        5'd0: x23y0 = in;
                        5'd1: x23y1 = in;
                        5'd2: x23y2 = in;
                        5'd3: x23y3 = in;
                        5'd4: x23y4 = in;
                        5'd5: x23y5 = in;
                        5'd6: x23y6 = in;
                        5'd7: x23y7 = in;
                        5'd8: x23y8 = in;
                        5'd9: x23y9 = in;
                        5'd10: x23y10 = in;
                        5'd11: x23y11 = in;
                        5'd12: x23y12 = in;
                        5'd13: x23y13 = in;
                        5'd14: x23y14 = in;
                        5'd15: x23y15 = in;
                        5'd16: x23y16 = in;
                        5'd17: x23y17 = in;
                        5'd18: x23y18 = in;
                        5'd19: x23y19 = in;
                        5'd20: x23y20 = in;
                        5'd21: x23y21 = in;
                        5'd22: x23y22 = in;
                        5'd23: x23y23 = in;
                        5'd24: x23y24 = in;
                        5'd25: x23y25 = in;
                        5'd26: x23y26 = in;
                        5'd27: x23y27 = in;
                        5'd28: x23y28 = in;
                        5'd29: x23y29 = in;
                        default: ;
                    endcase
                end
                6'd24: begin
                    case (y)
                        5'd0: x24y0 = in;
                        5'd1: x24y1 = in;
                        5'd2: x24y2 = in;
                        5'd3: x24y3 = in;
                        5'd4: x24y4 = in;
                        5'd5: x24y5 = in;
                        5'd6: x24y6 = in;
                        5'd7: x24y7 = in;
                        5'd8: x24y8 = in;
                        5'd9: x24y9 = in;
                        5'd10: x24y10 = in;
                        5'd11: x24y11 = in;
                        5'd12: x24y12 = in;
                        5'd13: x24y13 = in;
                        5'd14: x24y14 = in;
                        5'd15: x24y15 = in;
                        5'd16: x24y16 = in;
                        5'd17: x24y17 = in;
                        5'd18: x24y18 = in;
                        5'd19: x24y19 = in;
                        5'd20: x24y20 = in;
                        5'd21: x24y21 = in;
                        5'd22: x24y22 = in;
                        5'd23: x24y23 = in;
                        5'd24: x24y24 = in;
                        5'd25: x24y25 = in;
                        5'd26: x24y26 = in;
                        5'd27: x24y27 = in;
                        5'd28: x24y28 = in;
                        5'd29: x24y29 = in;
                        default: ;
                    endcase
                end
                6'd25: begin
                    case (y)
                        5'd0: x25y0 = in;
                        5'd1: x25y1 = in;
                        5'd2: x25y2 = in;
                        5'd3: x25y3 = in;
                        5'd4: x25y4 = in;
                        5'd5: x25y5 = in;
                        5'd6: x25y6 = in;
                        5'd7: x25y7 = in;
                        5'd8: x25y8 = in;
                        5'd9: x25y9 = in;
                        5'd10: x25y10 = in;
                        5'd11: x25y11 = in;
                        5'd12: x25y12 = in;
                        5'd13: x25y13 = in;
                        5'd14: x25y14 = in;
                        5'd15: x25y15 = in;
                        5'd16: x25y16 = in;
                        5'd17: x25y17 = in;
                        5'd18: x25y18 = in;
                        5'd19: x25y19 = in;
                        5'd20: x25y20 = in;
                        5'd21: x25y21 = in;
                        5'd22: x25y22 = in;
                        5'd23: x25y23 = in;
                        5'd24: x25y24 = in;
                        5'd25: x25y25 = in;
                        5'd26: x25y26 = in;
                        5'd27: x25y27 = in;
                        5'd28: x25y28 = in;
                        5'd29: x25y29 = in;
                        default: ;
                    endcase
                end
                6'd26: begin
                    case (y)
                        5'd0: x26y0 = in;
                        5'd1: x26y1 = in;
                        5'd2: x26y2 = in;
                        5'd3: x26y3 = in;
                        5'd4: x26y4 = in;
                        5'd5: x26y5 = in;
                        5'd6: x26y6 = in;
                        5'd7: x26y7 = in;
                        5'd8: x26y8 = in;
                        5'd9: x26y9 = in;
                        5'd10: x26y10 = in;
                        5'd11: x26y11 = in;
                        5'd12: x26y12 = in;
                        5'd13: x26y13 = in;
                        5'd14: x26y14 = in;
                        5'd15: x26y15 = in;
                        5'd16: x26y16 = in;
                        5'd17: x26y17 = in;
                        5'd18: x26y18 = in;
                        5'd19: x26y19 = in;
                        5'd20: x26y20 = in;
                        5'd21: x26y21 = in;
                        5'd22: x26y22 = in;
                        5'd23: x26y23 = in;
                        5'd24: x26y24 = in;
                        5'd25: x26y25 = in;
                        5'd26: x26y26 = in;
                        5'd27: x26y27 = in;
                        5'd28: x26y28 = in;
                        5'd29: x26y29 = in;
                        default: ;
                    endcase
                end
                6'd27: begin
                    case (y)
                        5'd0: x27y0 = in;
                        5'd1: x27y1 = in;
                        5'd2: x27y2 = in;
                        5'd3: x27y3 = in;
                        5'd4: x27y4 = in;
                        5'd5: x27y5 = in;
                        5'd6: x27y6 = in;
                        5'd7: x27y7 = in;
                        5'd8: x27y8 = in;
                        5'd9: x27y9 = in;
                        5'd10: x27y10 = in;
                        5'd11: x27y11 = in;
                        5'd12: x27y12 = in;
                        5'd13: x27y13 = in;
                        5'd14: x27y14 = in;
                        5'd15: x27y15 = in;
                        5'd16: x27y16 = in;
                        5'd17: x27y17 = in;
                        5'd18: x27y18 = in;
                        5'd19: x27y19 = in;
                        5'd20: x27y20 = in;
                        5'd21: x27y21 = in;
                        5'd22: x27y22 = in;
                        5'd23: x27y23 = in;
                        5'd24: x27y24 = in;
                        5'd25: x27y25 = in;
                        5'd26: x27y26 = in;
                        5'd27: x27y27 = in;
                        5'd28: x27y28 = in;
                        5'd29: x27y29 = in;
                        default: ;
                    endcase
                end
                6'd28: begin
                    case (y)
                        5'd0: x28y0 = in;
                        5'd1: x28y1 = in;
                        5'd2: x28y2 = in;
                        5'd3: x28y3 = in;
                        5'd4: x28y4 = in;
                        5'd5: x28y5 = in;
                        5'd6: x28y6 = in;
                        5'd7: x28y7 = in;
                        5'd8: x28y8 = in;
                        5'd9: x28y9 = in;
                        5'd10: x28y10 = in;
                        5'd11: x28y11 = in;
                        5'd12: x28y12 = in;
                        5'd13: x28y13 = in;
                        5'd14: x28y14 = in;
                        5'd15: x28y15 = in;
                        5'd16: x28y16 = in;
                        5'd17: x28y17 = in;
                        5'd18: x28y18 = in;
                        5'd19: x28y19 = in;
                        5'd20: x28y20 = in;
                        5'd21: x28y21 = in;
                        5'd22: x28y22 = in;
                        5'd23: x28y23 = in;
                        5'd24: x28y24 = in;
                        5'd25: x28y25 = in;
                        5'd26: x28y26 = in;
                        5'd27: x28y27 = in;
                        5'd28: x28y28 = in;
                        5'd29: x28y29 = in;
                        default: ;
                    endcase
                end
                6'd29: begin
                    case (y)
                        5'd0: x29y0 = in;
                        5'd1: x29y1 = in;
                        5'd2: x29y2 = in;
                        5'd3: x29y3 = in;
                        5'd4: x29y4 = in;
                        5'd5: x29y5 = in;
                        5'd6: x29y6 = in;
                        5'd7: x29y7 = in;
                        5'd8: x29y8 = in;
                        5'd9: x29y9 = in;
                        5'd10: x29y10 = in;
                        5'd11: x29y11 = in;
                        5'd12: x29y12 = in;
                        5'd13: x29y13 = in;
                        5'd14: x29y14 = in;
                        5'd15: x29y15 = in;
                        5'd16: x29y16 = in;
                        5'd17: x29y17 = in;
                        5'd18: x29y18 = in;
                        5'd19: x29y19 = in;
                        5'd20: x29y20 = in;
                        5'd21: x29y21 = in;
                        5'd22: x29y22 = in;
                        5'd23: x29y23 = in;
                        5'd24: x29y24 = in;
                        5'd25: x29y25 = in;
                        5'd26: x29y26 = in;
                        5'd27: x29y27 = in;
                        5'd28: x29y28 = in;
                        5'd29: x29y29 = in;
                        default: ;
                    endcase
                end
                6'd30: begin
                    case (y)
                        5'd0: x30y0 = in;
                        5'd1: x30y1 = in;
                        5'd2: x30y2 = in;
                        5'd3: x30y3 = in;
                        5'd4: x30y4 = in;
                        5'd5: x30y5 = in;
                        5'd6: x30y6 = in;
                        5'd7: x30y7 = in;
                        5'd8: x30y8 = in;
                        5'd9: x30y9 = in;
                        5'd10: x30y10 = in;
                        5'd11: x30y11 = in;
                        5'd12: x30y12 = in;
                        5'd13: x30y13 = in;
                        5'd14: x30y14 = in;
                        5'd15: x30y15 = in;
                        5'd16: x30y16 = in;
                        5'd17: x30y17 = in;
                        5'd18: x30y18 = in;
                        5'd19: x30y19 = in;
                        5'd20: x30y20 = in;
                        5'd21: x30y21 = in;
                        5'd22: x30y22 = in;
                        5'd23: x30y23 = in;
                        5'd24: x30y24 = in;
                        5'd25: x30y25 = in;
                        5'd26: x30y26 = in;
                        5'd27: x30y27 = in;
                        5'd28: x30y28 = in;
                        5'd29: x30y29 = in;
                        default: ;
                    endcase
                end
                6'd31: begin
                    case (y)
                        5'd0: x31y0 = in;
                        5'd1: x31y1 = in;
                        5'd2: x31y2 = in;
                        5'd3: x31y3 = in;
                        5'd4: x31y4 = in;
                        5'd5: x31y5 = in;
                        5'd6: x31y6 = in;
                        5'd7: x31y7 = in;
                        5'd8: x31y8 = in;
                        5'd9: x31y9 = in;
                        5'd10: x31y10 = in;
                        5'd11: x31y11 = in;
                        5'd12: x31y12 = in;
                        5'd13: x31y13 = in;
                        5'd14: x31y14 = in;
                        5'd15: x31y15 = in;
                        5'd16: x31y16 = in;
                        5'd17: x31y17 = in;
                        5'd18: x31y18 = in;
                        5'd19: x31y19 = in;
                        5'd20: x31y20 = in;
                        5'd21: x31y21 = in;
                        5'd22: x31y22 = in;
                        5'd23: x31y23 = in;
                        5'd24: x31y24 = in;
                        5'd25: x31y25 = in;
                        5'd26: x31y26 = in;
                        5'd27: x31y27 = in;
                        5'd28: x31y28 = in;
                        5'd29: x31y29 = in;
                        default: ;
                    endcase
                end
                6'd32: begin
                    case (y)
                        5'd0: x32y0 = in;
                        5'd1: x32y1 = in;
                        5'd2: x32y2 = in;
                        5'd3: x32y3 = in;
                        5'd4: x32y4 = in;
                        5'd5: x32y5 = in;
                        5'd6: x32y6 = in;
                        5'd7: x32y7 = in;
                        5'd8: x32y8 = in;
                        5'd9: x32y9 = in;
                        5'd10: x32y10 = in;
                        5'd11: x32y11 = in;
                        5'd12: x32y12 = in;
                        5'd13: x32y13 = in;
                        5'd14: x32y14 = in;
                        5'd15: x32y15 = in;
                        5'd16: x32y16 = in;
                        5'd17: x32y17 = in;
                        5'd18: x32y18 = in;
                        5'd19: x32y19 = in;
                        5'd20: x32y20 = in;
                        5'd21: x32y21 = in;
                        5'd22: x32y22 = in;
                        5'd23: x32y23 = in;
                        5'd24: x32y24 = in;
                        5'd25: x32y25 = in;
                        5'd26: x32y26 = in;
                        5'd27: x32y27 = in;
                        5'd28: x32y28 = in;
                        5'd29: x32y29 = in;
                        default: ;
                    endcase
                end
                6'd33: begin
                    case (y)
                        5'd0: x33y0 = in;
                        5'd1: x33y1 = in;
                        5'd2: x33y2 = in;
                        5'd3: x33y3 = in;
                        5'd4: x33y4 = in;
                        5'd5: x33y5 = in;
                        5'd6: x33y6 = in;
                        5'd7: x33y7 = in;
                        5'd8: x33y8 = in;
                        5'd9: x33y9 = in;
                        5'd10: x33y10 = in;
                        5'd11: x33y11 = in;
                        5'd12: x33y12 = in;
                        5'd13: x33y13 = in;
                        5'd14: x33y14 = in;
                        5'd15: x33y15 = in;
                        5'd16: x33y16 = in;
                        5'd17: x33y17 = in;
                        5'd18: x33y18 = in;
                        5'd19: x33y19 = in;
                        5'd20: x33y20 = in;
                        5'd21: x33y21 = in;
                        5'd22: x33y22 = in;
                        5'd23: x33y23 = in;
                        5'd24: x33y24 = in;
                        5'd25: x33y25 = in;
                        5'd26: x33y26 = in;
                        5'd27: x33y27 = in;
                        5'd28: x33y28 = in;
                        5'd29: x33y29 = in;
                        default: ;
                    endcase
                end
                6'd34: begin
                    case (y)
                        5'd0: x34y0 = in;
                        5'd1: x34y1 = in;
                        5'd2: x34y2 = in;
                        5'd3: x34y3 = in;
                        5'd4: x34y4 = in;
                        5'd5: x34y5 = in;
                        5'd6: x34y6 = in;
                        5'd7: x34y7 = in;
                        5'd8: x34y8 = in;
                        5'd9: x34y9 = in;
                        5'd10: x34y10 = in;
                        5'd11: x34y11 = in;
                        5'd12: x34y12 = in;
                        5'd13: x34y13 = in;
                        5'd14: x34y14 = in;
                        5'd15: x34y15 = in;
                        5'd16: x34y16 = in;
                        5'd17: x34y17 = in;
                        5'd18: x34y18 = in;
                        5'd19: x34y19 = in;
                        5'd20: x34y20 = in;
                        5'd21: x34y21 = in;
                        5'd22: x34y22 = in;
                        5'd23: x34y23 = in;
                        5'd24: x34y24 = in;
                        5'd25: x34y25 = in;
                        5'd26: x34y26 = in;
                        5'd27: x34y27 = in;
                        5'd28: x34y28 = in;
                        5'd29: x34y29 = in;
                        default: ;
                    endcase
                end
                6'd35: begin
                    case (y)
                        5'd0: x35y0 = in;
                        5'd1: x35y1 = in;
                        5'd2: x35y2 = in;
                        5'd3: x35y3 = in;
                        5'd4: x35y4 = in;
                        5'd5: x35y5 = in;
                        5'd6: x35y6 = in;
                        5'd7: x35y7 = in;
                        5'd8: x35y8 = in;
                        5'd9: x35y9 = in;
                        5'd10: x35y10 = in;
                        5'd11: x35y11 = in;
                        5'd12: x35y12 = in;
                        5'd13: x35y13 = in;
                        5'd14: x35y14 = in;
                        5'd15: x35y15 = in;
                        5'd16: x35y16 = in;
                        5'd17: x35y17 = in;
                        5'd18: x35y18 = in;
                        5'd19: x35y19 = in;
                        5'd20: x35y20 = in;
                        5'd21: x35y21 = in;
                        5'd22: x35y22 = in;
                        5'd23: x35y23 = in;
                        5'd24: x35y24 = in;
                        5'd25: x35y25 = in;
                        5'd26: x35y26 = in;
                        5'd27: x35y27 = in;
                        5'd28: x35y28 = in;
                        5'd29: x35y29 = in;
                        default: ;
                    endcase
                end
                6'd36: begin
                    case (y)
                        5'd0: x36y0 = in;
                        5'd1: x36y1 = in;
                        5'd2: x36y2 = in;
                        5'd3: x36y3 = in;
                        5'd4: x36y4 = in;
                        5'd5: x36y5 = in;
                        5'd6: x36y6 = in;
                        5'd7: x36y7 = in;
                        5'd8: x36y8 = in;
                        5'd9: x36y9 = in;
                        5'd10: x36y10 = in;
                        5'd11: x36y11 = in;
                        5'd12: x36y12 = in;
                        5'd13: x36y13 = in;
                        5'd14: x36y14 = in;
                        5'd15: x36y15 = in;
                        5'd16: x36y16 = in;
                        5'd17: x36y17 = in;
                        5'd18: x36y18 = in;
                        5'd19: x36y19 = in;
                        5'd20: x36y20 = in;
                        5'd21: x36y21 = in;
                        5'd22: x36y22 = in;
                        5'd23: x36y23 = in;
                        5'd24: x36y24 = in;
                        5'd25: x36y25 = in;
                        5'd26: x36y26 = in;
                        5'd27: x36y27 = in;
                        5'd28: x36y28 = in;
                        5'd29: x36y29 = in;
                        default: ;
                    endcase
                end
                6'd37: begin
                    case (y)
                        5'd0: x37y0 = in;
                        5'd1: x37y1 = in;
                        5'd2: x37y2 = in;
                        5'd3: x37y3 = in;
                        5'd4: x37y4 = in;
                        5'd5: x37y5 = in;
                        5'd6: x37y6 = in;
                        5'd7: x37y7 = in;
                        5'd8: x37y8 = in;
                        5'd9: x37y9 = in;
                        5'd10: x37y10 = in;
                        5'd11: x37y11 = in;
                        5'd12: x37y12 = in;
                        5'd13: x37y13 = in;
                        5'd14: x37y14 = in;
                        5'd15: x37y15 = in;
                        5'd16: x37y16 = in;
                        5'd17: x37y17 = in;
                        5'd18: x37y18 = in;
                        5'd19: x37y19 = in;
                        5'd20: x37y20 = in;
                        5'd21: x37y21 = in;
                        5'd22: x37y22 = in;
                        5'd23: x37y23 = in;
                        5'd24: x37y24 = in;
                        5'd25: x37y25 = in;
                        5'd26: x37y26 = in;
                        5'd27: x37y27 = in;
                        5'd28: x37y28 = in;
                        5'd29: x37y29 = in;
                        default: ;
                    endcase
                end
                6'd38: begin
                    case (y)
                        5'd0: x38y0 = in;
                        5'd1: x38y1 = in;
                        5'd2: x38y2 = in;
                        5'd3: x38y3 = in;
                        5'd4: x38y4 = in;
                        5'd5: x38y5 = in;
                        5'd6: x38y6 = in;
                        5'd7: x38y7 = in;
                        5'd8: x38y8 = in;
                        5'd9: x38y9 = in;
                        5'd10: x38y10 = in;
                        5'd11: x38y11 = in;
                        5'd12: x38y12 = in;
                        5'd13: x38y13 = in;
                        5'd14: x38y14 = in;
                        5'd15: x38y15 = in;
                        5'd16: x38y16 = in;
                        5'd17: x38y17 = in;
                        5'd18: x38y18 = in;
                        5'd19: x38y19 = in;
                        5'd20: x38y20 = in;
                        5'd21: x38y21 = in;
                        5'd22: x38y22 = in;
                        5'd23: x38y23 = in;
                        5'd24: x38y24 = in;
                        5'd25: x38y25 = in;
                        5'd26: x38y26 = in;
                        5'd27: x38y27 = in;
                        5'd28: x38y28 = in;
                        5'd29: x38y29 = in;
                        default: ;
                    endcase
                end
                6'd39: begin
                    case (y)
                        5'd0: x39y0 = in;
                        5'd1: x39y1 = in;
                        5'd2: x39y2 = in;
                        5'd3: x39y3 = in;
                        5'd4: x39y4 = in;
                        5'd5: x39y5 = in;
                        5'd6: x39y6 = in;
                        5'd7: x39y7 = in;
                        5'd8: x39y8 = in;
                        5'd9: x39y9 = in;
                        5'd10: x39y10 = in;
                        5'd11: x39y11 = in;
                        5'd12: x39y12 = in;
                        5'd13: x39y13 = in;
                        5'd14: x39y14 = in;
                        5'd15: x39y15 = in;
                        5'd16: x39y16 = in;
                        5'd17: x39y17 = in;
                        5'd18: x39y18 = in;
                        5'd19: x39y19 = in;
                        5'd20: x39y20 = in;
                        5'd21: x39y21 = in;
                        5'd22: x39y22 = in;
                        5'd23: x39y23 = in;
                        5'd24: x39y24 = in;
                        5'd25: x39y25 = in;
                        5'd26: x39y26 = in;
                        5'd27: x39y27 = in;
                        5'd28: x39y28 = in;
                        5'd29: x39y29 = in;
                        default: ;
                    endcase
                end
                default: ;
            endcase
        end // if 

        // Reading address values, make sure to read everytime
        case (x)
            6'd0: begin
                case (y)
                    5'd0: out = x0y0;
                    5'd1: out = x0y1;
                    5'd2: out = x0y2;
                    5'd3: out = x0y3;
                    5'd4: out = x0y4;
                    5'd5: out = x0y5;
                    5'd6: out = x0y6;
                    5'd7: out = x0y7;
                    5'd8: out = x0y8;
                    5'd9: out = x0y9;
                    5'd10: out = x0y10;
                    5'd11: out = x0y11;
                    5'd12: out = x0y12;
                    5'd13: out = x0y13;
                    5'd14: out = x0y14;
                    5'd15: out = x0y15;
                    5'd16: out = x0y16;
                    5'd17: out = x0y17;
                    5'd18: out = x0y18;
                    5'd19: out = x0y19;
                    5'd20: out = x0y20;
                    5'd21: out = x0y21;
                    5'd22: out = x0y22;
                    5'd23: out = x0y23;
                    5'd24: out = x0y24;
                    5'd25: out = x0y25;
                    5'd26: out = x0y26;
                    5'd27: out = x0y27;
                    5'd28: out = x0y28;
                    5'd29: out = x0y29;
                    default: out = 3'd0;
                endcase
            end
            6'd1: begin
                case (y)
                    5'd0: out = x1y0;
                    5'd1: out = x1y1;
                    5'd2: out = x1y2;
                    5'd3: out = x1y3;
                    5'd4: out = x1y4;
                    5'd5: out = x1y5;
                    5'd6: out = x1y6;
                    5'd7: out = x1y7;
                    5'd8: out = x1y8;
                    5'd9: out = x1y9;
                    5'd10: out = x1y10;
                    5'd11: out = x1y11;
                    5'd12: out = x1y12;
                    5'd13: out = x1y13;
                    5'd14: out = x1y14;
                    5'd15: out = x1y15;
                    5'd16: out = x1y16;
                    5'd17: out = x1y17;
                    5'd18: out = x1y18;
                    5'd19: out = x1y19;
                    5'd20: out = x1y20;
                    5'd21: out = x1y21;
                    5'd22: out = x1y22;
                    5'd23: out = x1y23;
                    5'd24: out = x1y24;
                    5'd25: out = x1y25;
                    5'd26: out = x1y26;
                    5'd27: out = x1y27;
                    5'd28: out = x1y28;
                    5'd29: out = x1y29;
                    default: out = 3'd0;
                endcase
            end
            6'd2: begin
                case (y)
                    5'd0: out = x2y0;
                    5'd1: out = x2y1;
                    5'd2: out = x2y2;
                    5'd3: out = x2y3;
                    5'd4: out = x2y4;
                    5'd5: out = x2y5;
                    5'd6: out = x2y6;
                    5'd7: out = x2y7;
                    5'd8: out = x2y8;
                    5'd9: out = x2y9;
                    5'd10: out = x2y10;
                    5'd11: out = x2y11;
                    5'd12: out = x2y12;
                    5'd13: out = x2y13;
                    5'd14: out = x2y14;
                    5'd15: out = x2y15;
                    5'd16: out = x2y16;
                    5'd17: out = x2y17;
                    5'd18: out = x2y18;
                    5'd19: out = x2y19;
                    5'd20: out = x2y20;
                    5'd21: out = x2y21;
                    5'd22: out = x2y22;
                    5'd23: out = x2y23;
                    5'd24: out = x2y24;
                    5'd25: out = x2y25;
                    5'd26: out = x2y26;
                    5'd27: out = x2y27;
                    5'd28: out = x2y28;
                    5'd29: out = x2y29;
                    default: out = 3'd0;
                endcase
            end
            6'd3: begin
                case (y)
                    5'd0: out = x3y0;
                    5'd1: out = x3y1;
                    5'd2: out = x3y2;
                    5'd3: out = x3y3;
                    5'd4: out = x3y4;
                    5'd5: out = x3y5;
                    5'd6: out = x3y6;
                    5'd7: out = x3y7;
                    5'd8: out = x3y8;
                    5'd9: out = x3y9;
                    5'd10: out = x3y10;
                    5'd11: out = x3y11;
                    5'd12: out = x3y12;
                    5'd13: out = x3y13;
                    5'd14: out = x3y14;
                    5'd15: out = x3y15;
                    5'd16: out = x3y16;
                    5'd17: out = x3y17;
                    5'd18: out = x3y18;
                    5'd19: out = x3y19;
                    5'd20: out = x3y20;
                    5'd21: out = x3y21;
                    5'd22: out = x3y22;
                    5'd23: out = x3y23;
                    5'd24: out = x3y24;
                    5'd25: out = x3y25;
                    5'd26: out = x3y26;
                    5'd27: out = x3y27;
                    5'd28: out = x3y28;
                    5'd29: out = x3y29;
                    default: out = 3'd0;
                endcase
            end
            6'd4: begin
                case (y)
                    5'd0: out = x4y0;
                    5'd1: out = x4y1;
                    5'd2: out = x4y2;
                    5'd3: out = x4y3;
                    5'd4: out = x4y4;
                    5'd5: out = x4y5;
                    5'd6: out = x4y6;
                    5'd7: out = x4y7;
                    5'd8: out = x4y8;
                    5'd9: out = x4y9;
                    5'd10: out = x4y10;
                    5'd11: out = x4y11;
                    5'd12: out = x4y12;
                    5'd13: out = x4y13;
                    5'd14: out = x4y14;
                    5'd15: out = x4y15;
                    5'd16: out = x4y16;
                    5'd17: out = x4y17;
                    5'd18: out = x4y18;
                    5'd19: out = x4y19;
                    5'd20: out = x4y20;
                    5'd21: out = x4y21;
                    5'd22: out = x4y22;
                    5'd23: out = x4y23;
                    5'd24: out = x4y24;
                    5'd25: out = x4y25;
                    5'd26: out = x4y26;
                    5'd27: out = x4y27;
                    5'd28: out = x4y28;
                    5'd29: out = x4y29;
                    default: out = 3'd0;
                endcase
            end
            6'd5: begin
                case (y)
                    5'd0: out = x5y0;
                    5'd1: out = x5y1;
                    5'd2: out = x5y2;
                    5'd3: out = x5y3;
                    5'd4: out = x5y4;
                    5'd5: out = x5y5;
                    5'd6: out = x5y6;
                    5'd7: out = x5y7;
                    5'd8: out = x5y8;
                    5'd9: out = x5y9;
                    5'd10: out = x5y10;
                    5'd11: out = x5y11;
                    5'd12: out = x5y12;
                    5'd13: out = x5y13;
                    5'd14: out = x5y14;
                    5'd15: out = x5y15;
                    5'd16: out = x5y16;
                    5'd17: out = x5y17;
                    5'd18: out = x5y18;
                    5'd19: out = x5y19;
                    5'd20: out = x5y20;
                    5'd21: out = x5y21;
                    5'd22: out = x5y22;
                    5'd23: out = x5y23;
                    5'd24: out = x5y24;
                    5'd25: out = x5y25;
                    5'd26: out = x5y26;
                    5'd27: out = x5y27;
                    5'd28: out = x5y28;
                    5'd29: out = x5y29;
                    default: out = 3'd0;
                endcase
            end
            6'd6: begin
                case (y)
                    5'd0: out = x6y0;
                    5'd1: out = x6y1;
                    5'd2: out = x6y2;
                    5'd3: out = x6y3;
                    5'd4: out = x6y4;
                    5'd5: out = x6y5;
                    5'd6: out = x6y6;
                    5'd7: out = x6y7;
                    5'd8: out = x6y8;
                    5'd9: out = x6y9;
                    5'd10: out = x6y10;
                    5'd11: out = x6y11;
                    5'd12: out = x6y12;
                    5'd13: out = x6y13;
                    5'd14: out = x6y14;
                    5'd15: out = x6y15;
                    5'd16: out = x6y16;
                    5'd17: out = x6y17;
                    5'd18: out = x6y18;
                    5'd19: out = x6y19;
                    5'd20: out = x6y20;
                    5'd21: out = x6y21;
                    5'd22: out = x6y22;
                    5'd23: out = x6y23;
                    5'd24: out = x6y24;
                    5'd25: out = x6y25;
                    5'd26: out = x6y26;
                    5'd27: out = x6y27;
                    5'd28: out = x6y28;
                    5'd29: out = x6y29;
                    default: out = 3'd0;
                endcase
            end
            6'd7: begin
                case (y)
                    5'd0: out = x7y0;
                    5'd1: out = x7y1;
                    5'd2: out = x7y2;
                    5'd3: out = x7y3;
                    5'd4: out = x7y4;
                    5'd5: out = x7y5;
                    5'd6: out = x7y6;
                    5'd7: out = x7y7;
                    5'd8: out = x7y8;
                    5'd9: out = x7y9;
                    5'd10: out = x7y10;
                    5'd11: out = x7y11;
                    5'd12: out = x7y12;
                    5'd13: out = x7y13;
                    5'd14: out = x7y14;
                    5'd15: out = x7y15;
                    5'd16: out = x7y16;
                    5'd17: out = x7y17;
                    5'd18: out = x7y18;
                    5'd19: out = x7y19;
                    5'd20: out = x7y20;
                    5'd21: out = x7y21;
                    5'd22: out = x7y22;
                    5'd23: out = x7y23;
                    5'd24: out = x7y24;
                    5'd25: out = x7y25;
                    5'd26: out = x7y26;
                    5'd27: out = x7y27;
                    5'd28: out = x7y28;
                    5'd29: out = x7y29;
                    default: out = 3'd0;
                endcase
            end
            6'd8: begin
                case (y)
                    5'd0: out = x8y0;
                    5'd1: out = x8y1;
                    5'd2: out = x8y2;
                    5'd3: out = x8y3;
                    5'd4: out = x8y4;
                    5'd5: out = x8y5;
                    5'd6: out = x8y6;
                    5'd7: out = x8y7;
                    5'd8: out = x8y8;
                    5'd9: out = x8y9;
                    5'd10: out = x8y10;
                    5'd11: out = x8y11;
                    5'd12: out = x8y12;
                    5'd13: out = x8y13;
                    5'd14: out = x8y14;
                    5'd15: out = x8y15;
                    5'd16: out = x8y16;
                    5'd17: out = x8y17;
                    5'd18: out = x8y18;
                    5'd19: out = x8y19;
                    5'd20: out = x8y20;
                    5'd21: out = x8y21;
                    5'd22: out = x8y22;
                    5'd23: out = x8y23;
                    5'd24: out = x8y24;
                    5'd25: out = x8y25;
                    5'd26: out = x8y26;
                    5'd27: out = x8y27;
                    5'd28: out = x8y28;
                    5'd29: out = x8y29;
                    default: out = 3'd0;
                endcase
            end
            6'd9: begin
                case (y)
                    5'd0: out = x9y0;
                    5'd1: out = x9y1;
                    5'd2: out = x9y2;
                    5'd3: out = x9y3;
                    5'd4: out = x9y4;
                    5'd5: out = x9y5;
                    5'd6: out = x9y6;
                    5'd7: out = x9y7;
                    5'd8: out = x9y8;
                    5'd9: out = x9y9;
                    5'd10: out = x9y10;
                    5'd11: out = x9y11;
                    5'd12: out = x9y12;
                    5'd13: out = x9y13;
                    5'd14: out = x9y14;
                    5'd15: out = x9y15;
                    5'd16: out = x9y16;
                    5'd17: out = x9y17;
                    5'd18: out = x9y18;
                    5'd19: out = x9y19;
                    5'd20: out = x9y20;
                    5'd21: out = x9y21;
                    5'd22: out = x9y22;
                    5'd23: out = x9y23;
                    5'd24: out = x9y24;
                    5'd25: out = x9y25;
                    5'd26: out = x9y26;
                    5'd27: out = x9y27;
                    5'd28: out = x9y28;
                    5'd29: out = x9y29;
                    default: out = 3'd0;
                endcase
            end
            6'd10: begin
                case (y)
                    5'd0: out = x10y0;
                    5'd1: out = x10y1;
                    5'd2: out = x10y2;
                    5'd3: out = x10y3;
                    5'd4: out = x10y4;
                    5'd5: out = x10y5;
                    5'd6: out = x10y6;
                    5'd7: out = x10y7;
                    5'd8: out = x10y8;
                    5'd9: out = x10y9;
                    5'd10: out = x10y10;
                    5'd11: out = x10y11;
                    5'd12: out = x10y12;
                    5'd13: out = x10y13;
                    5'd14: out = x10y14;
                    5'd15: out = x10y15;
                    5'd16: out = x10y16;
                    5'd17: out = x10y17;
                    5'd18: out = x10y18;
                    5'd19: out = x10y19;
                    5'd20: out = x10y20;
                    5'd21: out = x10y21;
                    5'd22: out = x10y22;
                    5'd23: out = x10y23;
                    5'd24: out = x10y24;
                    5'd25: out = x10y25;
                    5'd26: out = x10y26;
                    5'd27: out = x10y27;
                    5'd28: out = x10y28;
                    5'd29: out = x10y29;
                    default: out = 3'd0;
                endcase
            end
            6'd11: begin
                case (y)
                    5'd0: out = x11y0;
                    5'd1: out = x11y1;
                    5'd2: out = x11y2;
                    5'd3: out = x11y3;
                    5'd4: out = x11y4;
                    5'd5: out = x11y5;
                    5'd6: out = x11y6;
                    5'd7: out = x11y7;
                    5'd8: out = x11y8;
                    5'd9: out = x11y9;
                    5'd10: out = x11y10;
                    5'd11: out = x11y11;
                    5'd12: out = x11y12;
                    5'd13: out = x11y13;
                    5'd14: out = x11y14;
                    5'd15: out = x11y15;
                    5'd16: out = x11y16;
                    5'd17: out = x11y17;
                    5'd18: out = x11y18;
                    5'd19: out = x11y19;
                    5'd20: out = x11y20;
                    5'd21: out = x11y21;
                    5'd22: out = x11y22;
                    5'd23: out = x11y23;
                    5'd24: out = x11y24;
                    5'd25: out = x11y25;
                    5'd26: out = x11y26;
                    5'd27: out = x11y27;
                    5'd28: out = x11y28;
                    5'd29: out = x11y29;
                    default: out = 3'd0;
                endcase
            end
            6'd12: begin
                case (y)
                    5'd0: out = x12y0;
                    5'd1: out = x12y1;
                    5'd2: out = x12y2;
                    5'd3: out = x12y3;
                    5'd4: out = x12y4;
                    5'd5: out = x12y5;
                    5'd6: out = x12y6;
                    5'd7: out = x12y7;
                    5'd8: out = x12y8;
                    5'd9: out = x12y9;
                    5'd10: out = x12y10;
                    5'd11: out = x12y11;
                    5'd12: out = x12y12;
                    5'd13: out = x12y13;
                    5'd14: out = x12y14;
                    5'd15: out = x12y15;
                    5'd16: out = x12y16;
                    5'd17: out = x12y17;
                    5'd18: out = x12y18;
                    5'd19: out = x12y19;
                    5'd20: out = x12y20;
                    5'd21: out = x12y21;
                    5'd22: out = x12y22;
                    5'd23: out = x12y23;
                    5'd24: out = x12y24;
                    5'd25: out = x12y25;
                    5'd26: out = x12y26;
                    5'd27: out = x12y27;
                    5'd28: out = x12y28;
                    5'd29: out = x12y29;
                    default: out = 3'd0;
                endcase
            end
            6'd13: begin
                case (y)
                    5'd0: out = x13y0;
                    5'd1: out = x13y1;
                    5'd2: out = x13y2;
                    5'd3: out = x13y3;
                    5'd4: out = x13y4;
                    5'd5: out = x13y5;
                    5'd6: out = x13y6;
                    5'd7: out = x13y7;
                    5'd8: out = x13y8;
                    5'd9: out = x13y9;
                    5'd10: out = x13y10;
                    5'd11: out = x13y11;
                    5'd12: out = x13y12;
                    5'd13: out = x13y13;
                    5'd14: out = x13y14;
                    5'd15: out = x13y15;
                    5'd16: out = x13y16;
                    5'd17: out = x13y17;
                    5'd18: out = x13y18;
                    5'd19: out = x13y19;
                    5'd20: out = x13y20;
                    5'd21: out = x13y21;
                    5'd22: out = x13y22;
                    5'd23: out = x13y23;
                    5'd24: out = x13y24;
                    5'd25: out = x13y25;
                    5'd26: out = x13y26;
                    5'd27: out = x13y27;
                    5'd28: out = x13y28;
                    5'd29: out = x13y29;
                    default: out = 3'd0;
                endcase
            end
            6'd14: begin
                case (y)
                    5'd0: out = x14y0;
                    5'd1: out = x14y1;
                    5'd2: out = x14y2;
                    5'd3: out = x14y3;
                    5'd4: out = x14y4;
                    5'd5: out = x14y5;
                    5'd6: out = x14y6;
                    5'd7: out = x14y7;
                    5'd8: out = x14y8;
                    5'd9: out = x14y9;
                    5'd10: out = x14y10;
                    5'd11: out = x14y11;
                    5'd12: out = x14y12;
                    5'd13: out = x14y13;
                    5'd14: out = x14y14;
                    5'd15: out = x14y15;
                    5'd16: out = x14y16;
                    5'd17: out = x14y17;
                    5'd18: out = x14y18;
                    5'd19: out = x14y19;
                    5'd20: out = x14y20;
                    5'd21: out = x14y21;
                    5'd22: out = x14y22;
                    5'd23: out = x14y23;
                    5'd24: out = x14y24;
                    5'd25: out = x14y25;
                    5'd26: out = x14y26;
                    5'd27: out = x14y27;
                    5'd28: out = x14y28;
                    5'd29: out = x14y29;
                    default: out = 3'd0;
                endcase
            end
            6'd15: begin
                case (y)
                    5'd0: out = x15y0;
                    5'd1: out = x15y1;
                    5'd2: out = x15y2;
                    5'd3: out = x15y3;
                    5'd4: out = x15y4;
                    5'd5: out = x15y5;
                    5'd6: out = x15y6;
                    5'd7: out = x15y7;
                    5'd8: out = x15y8;
                    5'd9: out = x15y9;
                    5'd10: out = x15y10;
                    5'd11: out = x15y11;
                    5'd12: out = x15y12;
                    5'd13: out = x15y13;
                    5'd14: out = x15y14;
                    5'd15: out = x15y15;
                    5'd16: out = x15y16;
                    5'd17: out = x15y17;
                    5'd18: out = x15y18;
                    5'd19: out = x15y19;
                    5'd20: out = x15y20;
                    5'd21: out = x15y21;
                    5'd22: out = x15y22;
                    5'd23: out = x15y23;
                    5'd24: out = x15y24;
                    5'd25: out = x15y25;
                    5'd26: out = x15y26;
                    5'd27: out = x15y27;
                    5'd28: out = x15y28;
                    5'd29: out = x15y29;
                    default: out = 3'd0;
                endcase
            end
            6'd16: begin
                case (y)
                    5'd0: out = x16y0;
                    5'd1: out = x16y1;
                    5'd2: out = x16y2;
                    5'd3: out = x16y3;
                    5'd4: out = x16y4;
                    5'd5: out = x16y5;
                    5'd6: out = x16y6;
                    5'd7: out = x16y7;
                    5'd8: out = x16y8;
                    5'd9: out = x16y9;
                    5'd10: out = x16y10;
                    5'd11: out = x16y11;
                    5'd12: out = x16y12;
                    5'd13: out = x16y13;
                    5'd14: out = x16y14;
                    5'd15: out = x16y15;
                    5'd16: out = x16y16;
                    5'd17: out = x16y17;
                    5'd18: out = x16y18;
                    5'd19: out = x16y19;
                    5'd20: out = x16y20;
                    5'd21: out = x16y21;
                    5'd22: out = x16y22;
                    5'd23: out = x16y23;
                    5'd24: out = x16y24;
                    5'd25: out = x16y25;
                    5'd26: out = x16y26;
                    5'd27: out = x16y27;
                    5'd28: out = x16y28;
                    5'd29: out = x16y29;
                    default: out = 3'd0;
                endcase
            end
            6'd17: begin
                case (y)
                    5'd0: out = x17y0;
                    5'd1: out = x17y1;
                    5'd2: out = x17y2;
                    5'd3: out = x17y3;
                    5'd4: out = x17y4;
                    5'd5: out = x17y5;
                    5'd6: out = x17y6;
                    5'd7: out = x17y7;
                    5'd8: out = x17y8;
                    5'd9: out = x17y9;
                    5'd10: out = x17y10;
                    5'd11: out = x17y11;
                    5'd12: out = x17y12;
                    5'd13: out = x17y13;
                    5'd14: out = x17y14;
                    5'd15: out = x17y15;
                    5'd16: out = x17y16;
                    5'd17: out = x17y17;
                    5'd18: out = x17y18;
                    5'd19: out = x17y19;
                    5'd20: out = x17y20;
                    5'd21: out = x17y21;
                    5'd22: out = x17y22;
                    5'd23: out = x17y23;
                    5'd24: out = x17y24;
                    5'd25: out = x17y25;
                    5'd26: out = x17y26;
                    5'd27: out = x17y27;
                    5'd28: out = x17y28;
                    5'd29: out = x17y29;
                    default: out = 3'd0;
                endcase
            end
            6'd18: begin
                case (y)
                    5'd0: out = x18y0;
                    5'd1: out = x18y1;
                    5'd2: out = x18y2;
                    5'd3: out = x18y3;
                    5'd4: out = x18y4;
                    5'd5: out = x18y5;
                    5'd6: out = x18y6;
                    5'd7: out = x18y7;
                    5'd8: out = x18y8;
                    5'd9: out = x18y9;
                    5'd10: out = x18y10;
                    5'd11: out = x18y11;
                    5'd12: out = x18y12;
                    5'd13: out = x18y13;
                    5'd14: out = x18y14;
                    5'd15: out = x18y15;
                    5'd16: out = x18y16;
                    5'd17: out = x18y17;
                    5'd18: out = x18y18;
                    5'd19: out = x18y19;
                    5'd20: out = x18y20;
                    5'd21: out = x18y21;
                    5'd22: out = x18y22;
                    5'd23: out = x18y23;
                    5'd24: out = x18y24;
                    5'd25: out = x18y25;
                    5'd26: out = x18y26;
                    5'd27: out = x18y27;
                    5'd28: out = x18y28;
                    5'd29: out = x18y29;
                    default: out = 3'd0;
                endcase
            end
            6'd19: begin
                case (y)
                    5'd0: out = x19y0;
                    5'd1: out = x19y1;
                    5'd2: out = x19y2;
                    5'd3: out = x19y3;
                    5'd4: out = x19y4;
                    5'd5: out = x19y5;
                    5'd6: out = x19y6;
                    5'd7: out = x19y7;
                    5'd8: out = x19y8;
                    5'd9: out = x19y9;
                    5'd10: out = x19y10;
                    5'd11: out = x19y11;
                    5'd12: out = x19y12;
                    5'd13: out = x19y13;
                    5'd14: out = x19y14;
                    5'd15: out = x19y15;
                    5'd16: out = x19y16;
                    5'd17: out = x19y17;
                    5'd18: out = x19y18;
                    5'd19: out = x19y19;
                    5'd20: out = x19y20;
                    5'd21: out = x19y21;
                    5'd22: out = x19y22;
                    5'd23: out = x19y23;
                    5'd24: out = x19y24;
                    5'd25: out = x19y25;
                    5'd26: out = x19y26;
                    5'd27: out = x19y27;
                    5'd28: out = x19y28;
                    5'd29: out = x19y29;
                    default: out = 3'd0;
                endcase
            end
            6'd20: begin
                case (y)
                    5'd0: out = x20y0;
                    5'd1: out = x20y1;
                    5'd2: out = x20y2;
                    5'd3: out = x20y3;
                    5'd4: out = x20y4;
                    5'd5: out = x20y5;
                    5'd6: out = x20y6;
                    5'd7: out = x20y7;
                    5'd8: out = x20y8;
                    5'd9: out = x20y9;
                    5'd10: out = x20y10;
                    5'd11: out = x20y11;
                    5'd12: out = x20y12;
                    5'd13: out = x20y13;
                    5'd14: out = x20y14;
                    5'd15: out = x20y15;
                    5'd16: out = x20y16;
                    5'd17: out = x20y17;
                    5'd18: out = x20y18;
                    5'd19: out = x20y19;
                    5'd20: out = x20y20;
                    5'd21: out = x20y21;
                    5'd22: out = x20y22;
                    5'd23: out = x20y23;
                    5'd24: out = x20y24;
                    5'd25: out = x20y25;
                    5'd26: out = x20y26;
                    5'd27: out = x20y27;
                    5'd28: out = x20y28;
                    5'd29: out = x20y29;
                    default: out = 3'd0;
                endcase
            end
            6'd21: begin
                case (y)
                    5'd0: out = x21y0;
                    5'd1: out = x21y1;
                    5'd2: out = x21y2;
                    5'd3: out = x21y3;
                    5'd4: out = x21y4;
                    5'd5: out = x21y5;
                    5'd6: out = x21y6;
                    5'd7: out = x21y7;
                    5'd8: out = x21y8;
                    5'd9: out = x21y9;
                    5'd10: out = x21y10;
                    5'd11: out = x21y11;
                    5'd12: out = x21y12;
                    5'd13: out = x21y13;
                    5'd14: out = x21y14;
                    5'd15: out = x21y15;
                    5'd16: out = x21y16;
                    5'd17: out = x21y17;
                    5'd18: out = x21y18;
                    5'd19: out = x21y19;
                    5'd20: out = x21y20;
                    5'd21: out = x21y21;
                    5'd22: out = x21y22;
                    5'd23: out = x21y23;
                    5'd24: out = x21y24;
                    5'd25: out = x21y25;
                    5'd26: out = x21y26;
                    5'd27: out = x21y27;
                    5'd28: out = x21y28;
                    5'd29: out = x21y29;
                    default: out = 3'd0;
                endcase
            end
            6'd22: begin
                case (y)
                    5'd0: out = x22y0;
                    5'd1: out = x22y1;
                    5'd2: out = x22y2;
                    5'd3: out = x22y3;
                    5'd4: out = x22y4;
                    5'd5: out = x22y5;
                    5'd6: out = x22y6;
                    5'd7: out = x22y7;
                    5'd8: out = x22y8;
                    5'd9: out = x22y9;
                    5'd10: out = x22y10;
                    5'd11: out = x22y11;
                    5'd12: out = x22y12;
                    5'd13: out = x22y13;
                    5'd14: out = x22y14;
                    5'd15: out = x22y15;
                    5'd16: out = x22y16;
                    5'd17: out = x22y17;
                    5'd18: out = x22y18;
                    5'd19: out = x22y19;
                    5'd20: out = x22y20;
                    5'd21: out = x22y21;
                    5'd22: out = x22y22;
                    5'd23: out = x22y23;
                    5'd24: out = x22y24;
                    5'd25: out = x22y25;
                    5'd26: out = x22y26;
                    5'd27: out = x22y27;
                    5'd28: out = x22y28;
                    5'd29: out = x22y29;
                    default: out = 3'd0;
                endcase
            end
            6'd23: begin
                case (y)
                    5'd0: out = x23y0;
                    5'd1: out = x23y1;
                    5'd2: out = x23y2;
                    5'd3: out = x23y3;
                    5'd4: out = x23y4;
                    5'd5: out = x23y5;
                    5'd6: out = x23y6;
                    5'd7: out = x23y7;
                    5'd8: out = x23y8;
                    5'd9: out = x23y9;
                    5'd10: out = x23y10;
                    5'd11: out = x23y11;
                    5'd12: out = x23y12;
                    5'd13: out = x23y13;
                    5'd14: out = x23y14;
                    5'd15: out = x23y15;
                    5'd16: out = x23y16;
                    5'd17: out = x23y17;
                    5'd18: out = x23y18;
                    5'd19: out = x23y19;
                    5'd20: out = x23y20;
                    5'd21: out = x23y21;
                    5'd22: out = x23y22;
                    5'd23: out = x23y23;
                    5'd24: out = x23y24;
                    5'd25: out = x23y25;
                    5'd26: out = x23y26;
                    5'd27: out = x23y27;
                    5'd28: out = x23y28;
                    5'd29: out = x23y29;
                    default: out = 3'd0;
                endcase
            end
            6'd24: begin
                case (y)
                    5'd0: out = x24y0;
                    5'd1: out = x24y1;
                    5'd2: out = x24y2;
                    5'd3: out = x24y3;
                    5'd4: out = x24y4;
                    5'd5: out = x24y5;
                    5'd6: out = x24y6;
                    5'd7: out = x24y7;
                    5'd8: out = x24y8;
                    5'd9: out = x24y9;
                    5'd10: out = x24y10;
                    5'd11: out = x24y11;
                    5'd12: out = x24y12;
                    5'd13: out = x24y13;
                    5'd14: out = x24y14;
                    5'd15: out = x24y15;
                    5'd16: out = x24y16;
                    5'd17: out = x24y17;
                    5'd18: out = x24y18;
                    5'd19: out = x24y19;
                    5'd20: out = x24y20;
                    5'd21: out = x24y21;
                    5'd22: out = x24y22;
                    5'd23: out = x24y23;
                    5'd24: out = x24y24;
                    5'd25: out = x24y25;
                    5'd26: out = x24y26;
                    5'd27: out = x24y27;
                    5'd28: out = x24y28;
                    5'd29: out = x24y29;
                    default: out = 3'd0;
                endcase
            end
            6'd25: begin
                case (y)
                    5'd0: out = x25y0;
                    5'd1: out = x25y1;
                    5'd2: out = x25y2;
                    5'd3: out = x25y3;
                    5'd4: out = x25y4;
                    5'd5: out = x25y5;
                    5'd6: out = x25y6;
                    5'd7: out = x25y7;
                    5'd8: out = x25y8;
                    5'd9: out = x25y9;
                    5'd10: out = x25y10;
                    5'd11: out = x25y11;
                    5'd12: out = x25y12;
                    5'd13: out = x25y13;
                    5'd14: out = x25y14;
                    5'd15: out = x25y15;
                    5'd16: out = x25y16;
                    5'd17: out = x25y17;
                    5'd18: out = x25y18;
                    5'd19: out = x25y19;
                    5'd20: out = x25y20;
                    5'd21: out = x25y21;
                    5'd22: out = x25y22;
                    5'd23: out = x25y23;
                    5'd24: out = x25y24;
                    5'd25: out = x25y25;
                    5'd26: out = x25y26;
                    5'd27: out = x25y27;
                    5'd28: out = x25y28;
                    5'd29: out = x25y29;
                    default: out = 3'd0;
                endcase
            end
            6'd26: begin
                case (y)
                    5'd0: out = x26y0;
                    5'd1: out = x26y1;
                    5'd2: out = x26y2;
                    5'd3: out = x26y3;
                    5'd4: out = x26y4;
                    5'd5: out = x26y5;
                    5'd6: out = x26y6;
                    5'd7: out = x26y7;
                    5'd8: out = x26y8;
                    5'd9: out = x26y9;
                    5'd10: out = x26y10;
                    5'd11: out = x26y11;
                    5'd12: out = x26y12;
                    5'd13: out = x26y13;
                    5'd14: out = x26y14;
                    5'd15: out = x26y15;
                    5'd16: out = x26y16;
                    5'd17: out = x26y17;
                    5'd18: out = x26y18;
                    5'd19: out = x26y19;
                    5'd20: out = x26y20;
                    5'd21: out = x26y21;
                    5'd22: out = x26y22;
                    5'd23: out = x26y23;
                    5'd24: out = x26y24;
                    5'd25: out = x26y25;
                    5'd26: out = x26y26;
                    5'd27: out = x26y27;
                    5'd28: out = x26y28;
                    5'd29: out = x26y29;
                    default: out = 3'd0;
                endcase
            end
            6'd27: begin
                case (y)
                    5'd0: out = x27y0;
                    5'd1: out = x27y1;
                    5'd2: out = x27y2;
                    5'd3: out = x27y3;
                    5'd4: out = x27y4;
                    5'd5: out = x27y5;
                    5'd6: out = x27y6;
                    5'd7: out = x27y7;
                    5'd8: out = x27y8;
                    5'd9: out = x27y9;
                    5'd10: out = x27y10;
                    5'd11: out = x27y11;
                    5'd12: out = x27y12;
                    5'd13: out = x27y13;
                    5'd14: out = x27y14;
                    5'd15: out = x27y15;
                    5'd16: out = x27y16;
                    5'd17: out = x27y17;
                    5'd18: out = x27y18;
                    5'd19: out = x27y19;
                    5'd20: out = x27y20;
                    5'd21: out = x27y21;
                    5'd22: out = x27y22;
                    5'd23: out = x27y23;
                    5'd24: out = x27y24;
                    5'd25: out = x27y25;
                    5'd26: out = x27y26;
                    5'd27: out = x27y27;
                    5'd28: out = x27y28;
                    5'd29: out = x27y29;
                    default: out = 3'd0;
                endcase
            end
            6'd28: begin
                case (y)
                    5'd0: out = x28y0;
                    5'd1: out = x28y1;
                    5'd2: out = x28y2;
                    5'd3: out = x28y3;
                    5'd4: out = x28y4;
                    5'd5: out = x28y5;
                    5'd6: out = x28y6;
                    5'd7: out = x28y7;
                    5'd8: out = x28y8;
                    5'd9: out = x28y9;
                    5'd10: out = x28y10;
                    5'd11: out = x28y11;
                    5'd12: out = x28y12;
                    5'd13: out = x28y13;
                    5'd14: out = x28y14;
                    5'd15: out = x28y15;
                    5'd16: out = x28y16;
                    5'd17: out = x28y17;
                    5'd18: out = x28y18;
                    5'd19: out = x28y19;
                    5'd20: out = x28y20;
                    5'd21: out = x28y21;
                    5'd22: out = x28y22;
                    5'd23: out = x28y23;
                    5'd24: out = x28y24;
                    5'd25: out = x28y25;
                    5'd26: out = x28y26;
                    5'd27: out = x28y27;
                    5'd28: out = x28y28;
                    5'd29: out = x28y29;
                    default: out = 3'd0;
                endcase
            end
            6'd29: begin
                case (y)
                    5'd0: out = x29y0;
                    5'd1: out = x29y1;
                    5'd2: out = x29y2;
                    5'd3: out = x29y3;
                    5'd4: out = x29y4;
                    5'd5: out = x29y5;
                    5'd6: out = x29y6;
                    5'd7: out = x29y7;
                    5'd8: out = x29y8;
                    5'd9: out = x29y9;
                    5'd10: out = x29y10;
                    5'd11: out = x29y11;
                    5'd12: out = x29y12;
                    5'd13: out = x29y13;
                    5'd14: out = x29y14;
                    5'd15: out = x29y15;
                    5'd16: out = x29y16;
                    5'd17: out = x29y17;
                    5'd18: out = x29y18;
                    5'd19: out = x29y19;
                    5'd20: out = x29y20;
                    5'd21: out = x29y21;
                    5'd22: out = x29y22;
                    5'd23: out = x29y23;
                    5'd24: out = x29y24;
                    5'd25: out = x29y25;
                    5'd26: out = x29y26;
                    5'd27: out = x29y27;
                    5'd28: out = x29y28;
                    5'd29: out = x29y29;
                    default: out = 3'd0;
                endcase
            end
            6'd30: begin
                case (y)
                    5'd0: out = x30y0;
                    5'd1: out = x30y1;
                    5'd2: out = x30y2;
                    5'd3: out = x30y3;
                    5'd4: out = x30y4;
                    5'd5: out = x30y5;
                    5'd6: out = x30y6;
                    5'd7: out = x30y7;
                    5'd8: out = x30y8;
                    5'd9: out = x30y9;
                    5'd10: out = x30y10;
                    5'd11: out = x30y11;
                    5'd12: out = x30y12;
                    5'd13: out = x30y13;
                    5'd14: out = x30y14;
                    5'd15: out = x30y15;
                    5'd16: out = x30y16;
                    5'd17: out = x30y17;
                    5'd18: out = x30y18;
                    5'd19: out = x30y19;
                    5'd20: out = x30y20;
                    5'd21: out = x30y21;
                    5'd22: out = x30y22;
                    5'd23: out = x30y23;
                    5'd24: out = x30y24;
                    5'd25: out = x30y25;
                    5'd26: out = x30y26;
                    5'd27: out = x30y27;
                    5'd28: out = x30y28;
                    5'd29: out = x30y29;
                    default: out = 3'd0;
                endcase
            end
            6'd31: begin
                case (y)
                    5'd0: out = x31y0;
                    5'd1: out = x31y1;
                    5'd2: out = x31y2;
                    5'd3: out = x31y3;
                    5'd4: out = x31y4;
                    5'd5: out = x31y5;
                    5'd6: out = x31y6;
                    5'd7: out = x31y7;
                    5'd8: out = x31y8;
                    5'd9: out = x31y9;
                    5'd10: out = x31y10;
                    5'd11: out = x31y11;
                    5'd12: out = x31y12;
                    5'd13: out = x31y13;
                    5'd14: out = x31y14;
                    5'd15: out = x31y15;
                    5'd16: out = x31y16;
                    5'd17: out = x31y17;
                    5'd18: out = x31y18;
                    5'd19: out = x31y19;
                    5'd20: out = x31y20;
                    5'd21: out = x31y21;
                    5'd22: out = x31y22;
                    5'd23: out = x31y23;
                    5'd24: out = x31y24;
                    5'd25: out = x31y25;
                    5'd26: out = x31y26;
                    5'd27: out = x31y27;
                    5'd28: out = x31y28;
                    5'd29: out = x31y29;
                    default: out = 3'd0;
                endcase
            end
            6'd32: begin
                case (y)
                    5'd0: out = x32y0;
                    5'd1: out = x32y1;
                    5'd2: out = x32y2;
                    5'd3: out = x32y3;
                    5'd4: out = x32y4;
                    5'd5: out = x32y5;
                    5'd6: out = x32y6;
                    5'd7: out = x32y7;
                    5'd8: out = x32y8;
                    5'd9: out = x32y9;
                    5'd10: out = x32y10;
                    5'd11: out = x32y11;
                    5'd12: out = x32y12;
                    5'd13: out = x32y13;
                    5'd14: out = x32y14;
                    5'd15: out = x32y15;
                    5'd16: out = x32y16;
                    5'd17: out = x32y17;
                    5'd18: out = x32y18;
                    5'd19: out = x32y19;
                    5'd20: out = x32y20;
                    5'd21: out = x32y21;
                    5'd22: out = x32y22;
                    5'd23: out = x32y23;
                    5'd24: out = x32y24;
                    5'd25: out = x32y25;
                    5'd26: out = x32y26;
                    5'd27: out = x32y27;
                    5'd28: out = x32y28;
                    5'd29: out = x32y29;
                    default: out = 3'd0;
                endcase
            end
            6'd33: begin
                case (y)
                    5'd0: out = x33y0;
                    5'd1: out = x33y1;
                    5'd2: out = x33y2;
                    5'd3: out = x33y3;
                    5'd4: out = x33y4;
                    5'd5: out = x33y5;
                    5'd6: out = x33y6;
                    5'd7: out = x33y7;
                    5'd8: out = x33y8;
                    5'd9: out = x33y9;
                    5'd10: out = x33y10;
                    5'd11: out = x33y11;
                    5'd12: out = x33y12;
                    5'd13: out = x33y13;
                    5'd14: out = x33y14;
                    5'd15: out = x33y15;
                    5'd16: out = x33y16;
                    5'd17: out = x33y17;
                    5'd18: out = x33y18;
                    5'd19: out = x33y19;
                    5'd20: out = x33y20;
                    5'd21: out = x33y21;
                    5'd22: out = x33y22;
                    5'd23: out = x33y23;
                    5'd24: out = x33y24;
                    5'd25: out = x33y25;
                    5'd26: out = x33y26;
                    5'd27: out = x33y27;
                    5'd28: out = x33y28;
                    5'd29: out = x33y29;
                    default: out = 3'd0;
                endcase
            end
            6'd34: begin
                case (y)
                    5'd0: out = x34y0;
                    5'd1: out = x34y1;
                    5'd2: out = x34y2;
                    5'd3: out = x34y3;
                    5'd4: out = x34y4;
                    5'd5: out = x34y5;
                    5'd6: out = x34y6;
                    5'd7: out = x34y7;
                    5'd8: out = x34y8;
                    5'd9: out = x34y9;
                    5'd10: out = x34y10;
                    5'd11: out = x34y11;
                    5'd12: out = x34y12;
                    5'd13: out = x34y13;
                    5'd14: out = x34y14;
                    5'd15: out = x34y15;
                    5'd16: out = x34y16;
                    5'd17: out = x34y17;
                    5'd18: out = x34y18;
                    5'd19: out = x34y19;
                    5'd20: out = x34y20;
                    5'd21: out = x34y21;
                    5'd22: out = x34y22;
                    5'd23: out = x34y23;
                    5'd24: out = x34y24;
                    5'd25: out = x34y25;
                    5'd26: out = x34y26;
                    5'd27: out = x34y27;
                    5'd28: out = x34y28;
                    5'd29: out = x34y29;
                    default: out = 3'd0;
                endcase
            end
            6'd35: begin
                case (y)
                    5'd0: out = x35y0;
                    5'd1: out = x35y1;
                    5'd2: out = x35y2;
                    5'd3: out = x35y3;
                    5'd4: out = x35y4;
                    5'd5: out = x35y5;
                    5'd6: out = x35y6;
                    5'd7: out = x35y7;
                    5'd8: out = x35y8;
                    5'd9: out = x35y9;
                    5'd10: out = x35y10;
                    5'd11: out = x35y11;
                    5'd12: out = x35y12;
                    5'd13: out = x35y13;
                    5'd14: out = x35y14;
                    5'd15: out = x35y15;
                    5'd16: out = x35y16;
                    5'd17: out = x35y17;
                    5'd18: out = x35y18;
                    5'd19: out = x35y19;
                    5'd20: out = x35y20;
                    5'd21: out = x35y21;
                    5'd22: out = x35y22;
                    5'd23: out = x35y23;
                    5'd24: out = x35y24;
                    5'd25: out = x35y25;
                    5'd26: out = x35y26;
                    5'd27: out = x35y27;
                    5'd28: out = x35y28;
                    5'd29: out = x35y29;
                    default: out = 3'd0;
                endcase
            end
            6'd36: begin
                case (y)
                    5'd0: out = x36y0;
                    5'd1: out = x36y1;
                    5'd2: out = x36y2;
                    5'd3: out = x36y3;
                    5'd4: out = x36y4;
                    5'd5: out = x36y5;
                    5'd6: out = x36y6;
                    5'd7: out = x36y7;
                    5'd8: out = x36y8;
                    5'd9: out = x36y9;
                    5'd10: out = x36y10;
                    5'd11: out = x36y11;
                    5'd12: out = x36y12;
                    5'd13: out = x36y13;
                    5'd14: out = x36y14;
                    5'd15: out = x36y15;
                    5'd16: out = x36y16;
                    5'd17: out = x36y17;
                    5'd18: out = x36y18;
                    5'd19: out = x36y19;
                    5'd20: out = x36y20;
                    5'd21: out = x36y21;
                    5'd22: out = x36y22;
                    5'd23: out = x36y23;
                    5'd24: out = x36y24;
                    5'd25: out = x36y25;
                    5'd26: out = x36y26;
                    5'd27: out = x36y27;
                    5'd28: out = x36y28;
                    5'd29: out = x36y29;
                    default: out = 3'd0;
                endcase
            end
            6'd37: begin
                case (y)
                    5'd0: out = x37y0;
                    5'd1: out = x37y1;
                    5'd2: out = x37y2;
                    5'd3: out = x37y3;
                    5'd4: out = x37y4;
                    5'd5: out = x37y5;
                    5'd6: out = x37y6;
                    5'd7: out = x37y7;
                    5'd8: out = x37y8;
                    5'd9: out = x37y9;
                    5'd10: out = x37y10;
                    5'd11: out = x37y11;
                    5'd12: out = x37y12;
                    5'd13: out = x37y13;
                    5'd14: out = x37y14;
                    5'd15: out = x37y15;
                    5'd16: out = x37y16;
                    5'd17: out = x37y17;
                    5'd18: out = x37y18;
                    5'd19: out = x37y19;
                    5'd20: out = x37y20;
                    5'd21: out = x37y21;
                    5'd22: out = x37y22;
                    5'd23: out = x37y23;
                    5'd24: out = x37y24;
                    5'd25: out = x37y25;
                    5'd26: out = x37y26;
                    5'd27: out = x37y27;
                    5'd28: out = x37y28;
                    5'd29: out = x37y29;
                    default: out = 3'd0;
                endcase
            end
            6'd38: begin
                case (y)
                    5'd0: out = x38y0;
                    5'd1: out = x38y1;
                    5'd2: out = x38y2;
                    5'd3: out = x38y3;
                    5'd4: out = x38y4;
                    5'd5: out = x38y5;
                    5'd6: out = x38y6;
                    5'd7: out = x38y7;
                    5'd8: out = x38y8;
                    5'd9: out = x38y9;
                    5'd10: out = x38y10;
                    5'd11: out = x38y11;
                    5'd12: out = x38y12;
                    5'd13: out = x38y13;
                    5'd14: out = x38y14;
                    5'd15: out = x38y15;
                    5'd16: out = x38y16;
                    5'd17: out = x38y17;
                    5'd18: out = x38y18;
                    5'd19: out = x38y19;
                    5'd20: out = x38y20;
                    5'd21: out = x38y21;
                    5'd22: out = x38y22;
                    5'd23: out = x38y23;
                    5'd24: out = x38y24;
                    5'd25: out = x38y25;
                    5'd26: out = x38y26;
                    5'd27: out = x38y27;
                    5'd28: out = x38y28;
                    5'd29: out = x38y29;
                    default: out = 3'd0;
                endcase
            end
            6'd39: begin
                case (y)
                    5'd0: out = x39y0;
                    5'd1: out = x39y1;
                    5'd2: out = x39y2;
                    5'd3: out = x39y3;
                    5'd4: out = x39y4;
                    5'd5: out = x39y5;
                    5'd6: out = x39y6;
                    5'd7: out = x39y7;
                    5'd8: out = x39y8;
                    5'd9: out = x39y9;
                    5'd10: out = x39y10;
                    5'd11: out = x39y11;
                    5'd12: out = x39y12;
                    5'd13: out = x39y13;
                    5'd14: out = x39y14;
                    5'd15: out = x39y15;
                    5'd16: out = x39y16;
                    5'd17: out = x39y17;
                    5'd18: out = x39y18;
                    5'd19: out = x39y19;
                    5'd20: out = x39y20;
                    5'd21: out = x39y21;
                    5'd22: out = x39y22;
                    5'd23: out = x39y23;
                    5'd24: out = x39y24;
                    5'd25: out = x39y25;
                    5'd26: out = x39y26;
                    5'd27: out = x39y27;
                    5'd28: out = x39y28;
                    5'd29: out = x39y29;
                    default: out = 3'd0;
                endcase
            end
            default: out = 3'd0;
        endcase
    end // always
endmodule
