module player_updater(clock, reset,
                      start, done,
                      cur_pos_x, cur_pos_y, cur_angle,
                      next_pos_x, next_pos_y, next_angle,
                      grid_x, grid_y, grid_out);
    input clock;
    input reset;

    // Current player position and angle
    input [13:0] cur_pos_x;
    input [12:0] cur_pos_y;
    input [7:0] cur_angle;

    // Next player position and angle
    output [13:0] next_pos_x;
    output [12:0] next_pos_y;
    output [7:0] next_angle;

    output [5:0] grid_x;
    output [4:0] grid_y;
    input [2:0] grid_out;

    // TODO: Keyboard inputs
endmodule
