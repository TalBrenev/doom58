module level_loader(clock, start, level, grid_x, grid_y, grid_in, grid_write, done);
endmodule
