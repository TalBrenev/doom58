module level_loader(clock, reset, start, level, grid_x, grid_y, grid_in, grid_write, done);
endmodule
