module draw_grid(clock, start, grid_x, grid_y, grid_write, grid_out, vga_x, vga_y, vga_colour, vga_write, done);
endmodule
