module raytracer(clock, reset,
                 start, done,
                 x, y, angle,
                 grid_x, grid_y, grid_out);
endmodule
