module grid(clock, reset, x, y, write, in, out);
endmodule
