module grid(clock, x, y, write, in, out);
endmodule
