module raytracer(clock, start, x, y, angle, grid_x, grid_y, grid_write, grid_out, done);
endmodule
