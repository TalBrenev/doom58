module level_loader(clock, reset,
                    start, done,
                    level,
                    grid_x, grid_y, grid_in, grid_write);
endmodule
