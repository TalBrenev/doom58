module bytian_to_vector(bytian, x, y);
    input [7:0] bytian;

    output [13:0] x;
    output [12:0] y;
endmodule
